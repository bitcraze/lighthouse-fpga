module chip (io_12_31_1, io_13_31_0, io_17_0_0, io_17_31_0, io_18_0_0, io_18_31_1, io_22_0_1, io_6_0_0, io_7_0_0, io_8_31_1);
  wire net_5;
  wire net_6;
  wire net_8;
  wire net_10;
  wire net_11;
  wire net_1816;
  wire net_2864;
  wire net_7745;
  wire net_7746;
  wire net_7747;
  wire net_7748;
  wire net_7749;
  wire net_7750;
  wire net_9360;
  wire net_11035;
  wire net_11052;
  wire net_12015;
  wire net_12035;
  wire net_12039;
  wire net_12135;
  wire net_12178;
  wire net_12179;
  wire net_12185;
  wire net_12191;
  wire net_12192;
  wire net_12198;
  wire net_12200;
  wire net_12201;
  wire net_12206;
  wire net_12210;
  wire net_12213;
  wire net_12216;
  wire net_12218;
  wire net_12220;
  wire net_12222;
  wire net_12225;
  wire net_12226;
  wire net_12228;
  wire net_12231;
  wire net_12232;
  wire net_12236;
  wire net_12238;
  wire net_12241;
  wire net_12242;
  wire net_12243;
  wire net_12244;
  wire net_12247;
  wire net_12248;
  wire net_12249;
  wire net_12252;
  wire net_12253;
  wire net_12748;
  wire net_12749;
  wire net_12750;
  wire net_12751;
  wire net_12752;
  wire net_12753;
  wire net_12871;
  wire net_12886;
  wire net_13363;
  wire net_13364;
  wire net_13365;
  wire net_13366;
  wire net_13367;
  wire net_13368;
  wire net_13484;
  wire net_13485;
  wire net_13486;
  wire net_13487;
  wire net_13488;
  wire net_13489;
  wire net_13490;
  wire net_13491;
  wire net_13545;
  wire net_13551;
  wire net_13554;
  wire net_13555;
  wire net_13558;
  wire net_13559;
  wire net_13560;
  wire net_13561;
  wire net_13607;
  wire net_13608;
  wire net_13609;
  wire net_13610;
  wire net_13611;
  wire net_13612;
  wire net_13613;
  wire net_13614;
  wire net_13619;
  wire net_15887;
  wire net_15893;
  wire net_15895;
  wire net_15955;
  wire net_15958;
  wire net_15960;
  wire net_15961;
  wire net_16014;
  wire net_16015;
  wire net_16016;
  wire net_16061;
  wire net_16082;
  wire net_16083;
  wire net_16084;
  wire net_16095;
  wire net_16366;
  wire net_16456;
  wire net_16582;
  wire net_16620;
  wire net_16628;
  wire net_16631;
  wire net_16632;
  wire net_16639;
  wire net_16645;
  wire net_16646;
  wire net_16647;
  wire net_16652;
  wire net_16656;
  wire net_16659;
  wire net_16662;
  wire net_16665;
  wire net_16666;
  wire net_16668;
  wire net_16670;
  wire net_16672;
  wire net_16674;
  wire net_16676;
  wire net_16678;
  wire net_16682;
  wire net_16684;
  wire net_16687;
  wire net_16688;
  wire net_16689;
  wire net_16690;
  wire net_16693;
  wire net_16694;
  wire net_16695;
  wire net_16698;
  wire net_16699;
  wire net_16759;
  wire net_16768;
  wire net_16770;
  wire net_16786;
  wire net_16820;
  wire net_16821;
  wire net_16822;
  wire net_17070;
  wire net_17095;
  wire net_17192;
  wire net_17194;
  wire net_17198;
  wire net_17199;
  wire net_17237;
  wire net_17238;
  wire net_17239;
  wire net_17242;
  wire net_17251;
  wire net_17252;
  wire net_17256;
  wire net_17264;
  wire net_17267;
  wire net_17271;
  wire net_17273;
  wire net_17277;
  wire net_17280;
  wire net_17281;
  wire net_17283;
  wire net_17286;
  wire net_17287;
  wire net_17289;
  wire net_17292;
  wire net_17293;
  wire net_17295;
  wire net_17298;
  wire net_17299;
  wire net_17301;
  wire net_17304;
  wire net_17305;
  wire net_17307;
  wire net_17309;
  wire net_17311;
  wire net_17313;
  wire net_17316;
  wire net_17317;
  wire net_17319;
  wire net_17351;
  wire net_17357;
  wire net_17362;
  wire net_17364;
  wire net_17367;
  wire net_17376;
  wire net_17377;
  wire net_17379;
  wire net_17382;
  wire net_17388;
  wire net_17390;
  wire net_17392;
  wire net_17394;
  wire net_17397;
  wire net_17398;
  wire net_17400;
  wire net_17402;
  wire net_17404;
  wire net_17406;
  wire net_17408;
  wire net_17410;
  wire net_17412;
  wire net_17415;
  wire net_17416;
  wire net_17418;
  wire net_17421;
  wire net_17422;
  wire net_17424;
  wire net_17427;
  wire net_17428;
  wire net_17430;
  wire net_17433;
  wire net_17434;
  wire net_17436;
  wire net_17439;
  wire net_17474;
  wire net_17481;
  wire net_17493;
  wire net_17495;
  wire net_17500;
  wire net_17504;
  wire net_17506;
  wire net_17507;
  wire net_17510;
  wire net_17511;
  wire net_17514;
  wire net_17515;
  wire net_17517;
  wire net_17519;
  wire net_17521;
  wire net_17523;
  wire net_17526;
  wire net_17527;
  wire net_17529;
  wire net_17531;
  wire net_17533;
  wire net_17535;
  wire net_17537;
  wire net_17539;
  wire net_17541;
  wire net_17544;
  wire net_17545;
  wire net_17547;
  wire net_17549;
  wire net_17551;
  wire net_17555;
  wire net_17557;
  wire net_17559;
  wire net_19424;
  wire net_20287;
  wire net_20341;
  wire net_20352;
  wire net_20371;
  wire net_20374;
  wire net_20406;
  wire net_20426;
  wire net_20461;
  wire net_20462;
  wire net_20478;
  wire net_20513;
  wire net_20514;
  wire net_20529;
  wire net_20530;
  wire net_20805;
  wire net_20933;
  wire net_20942;
  wire net_20968;
  wire net_20982;
  wire net_21020;
  wire net_21021;
  wire net_21065;
  wire net_21066;
  wire net_21069;
  wire net_21070;
  wire net_21072;
  wire net_21073;
  wire net_21075;
  wire net_21076;
  wire net_21078;
  wire net_21086;
  wire net_21087;
  wire net_21089;
  wire net_21097;
  wire net_21098;
  wire net_21099;
  wire net_21100;
  wire net_21109;
  wire net_21111;
  wire net_21112;
  wire net_21133;
  wire net_21134;
  wire net_21135;
  wire net_21136;
  wire net_21139;
  wire net_21141;
  wire net_21144;
  wire net_21164;
  wire net_21171;
  wire net_21189;
  wire net_21190;
  wire net_21195;
  wire net_21196;
  wire net_21197;
  wire net_21199;
  wire net_21202;
  wire net_21203;
  wire net_21210;
  wire net_21211;
  wire net_21216;
  wire net_21218;
  wire net_21226;
  wire net_21227;
  wire net_21228;
  wire net_21229;
  wire net_21232;
  wire net_21233;
  wire net_21234;
  wire net_21235;
  wire net_21244;
  wire net_21245;
  wire net_21246;
  wire net_21247;
  wire net_21271;
  wire net_21313;
  wire net_21316;
  wire net_21319;
  wire net_21322;
  wire net_21349;
  wire net_21350;
  wire net_21351;
  wire net_21352;
  wire net_21400;
  wire net_22846;
  wire net_22847;
  wire net_22900;
  wire net_23161;
  wire net_23327;
  wire net_23331;
  wire net_23376;
  wire net_23390;
  wire net_24008;
  wire net_24159;
  wire net_24175;
  wire net_24202;
  wire net_24236;
  wire net_24237;
  wire net_24257;
  wire net_25152;
  wire net_25188;
  wire net_25220;
  wire net_25221;
  wire net_25241;
  wire net_26528;
  wire net_26534;
  wire net_26535;
  wire net_26536;
  wire net_26539;
  wire net_26547;
  wire net_26554;
  wire net_26571;
  wire net_26625;
  wire net_26691;
  wire net_26813;
  wire net_26919;
  wire net_27015;
  wire net_27633;
  wire net_27687;
  wire net_27688;
  wire net_27690;
  wire net_28343;
  wire net_29568;
  wire net_29728;
  wire net_29734;
  wire net_29735;
  wire net_29736;
  wire net_29743;
  wire net_29747;
  wire net_29814;
  wire net_29826;
  wire net_29836;
  wire net_29837;
  wire net_29882;
  wire net_29883;
  wire net_29884;
  wire net_29885;
  wire net_29886;
  wire net_29887;
  wire net_29888;
  wire net_29936;
  wire net_30041;
  wire net_30044;
  wire net_30045;
  wire net_30046;
  wire net_30047;
  wire net_30057;
  wire net_30164;
  wire net_30184;
  wire net_30198;
  wire net_30307;
  wire net_30790;
  wire net_30903;
  wire net_30904;
  wire net_30905;
  wire net_30906;
  wire net_30907;
  wire net_30908;
  wire net_30928;
  wire net_31029;
  wire net_31037;
  wire net_31041;
  wire net_31148;
  wire net_31207;
  wire net_31208;
  wire net_31213;
  wire net_31214;
  wire net_31223;
  wire net_31226;
  wire net_31228;
  wire net_31232;
  wire net_31234;
  wire net_31236;
  wire net_31239;
  wire net_31242;
  wire net_31251;
  wire net_31252;
  wire net_31253;
  wire net_31254;
  wire net_31268;
  wire net_31284;
  wire net_31767;
  wire net_32505;
  wire net_32527;
  wire net_32629;
  wire net_32748;
  wire net_32749;
  wire net_32750;
  wire net_32751;
  wire net_32752;
  wire net_32753;
  wire net_32775;
  wire net_32882;
  wire net_32901;
  wire net_33252;
  wire net_33486;
  wire net_33556;
  wire net_33712;
  wire net_33713;
  wire net_33714;
  wire net_33715;
  wire net_33716;
  wire net_33717;
  wire net_33718;
  wire net_33719;
  wire net_33722;
  wire net_33768;
  wire net_33774;
  wire net_33791;
  wire net_33797;
  wire net_33802;
  wire net_33803;
  wire net_33805;
  wire net_33814;
  wire net_33815;
  wire net_33816;
  wire net_33817;
  wire net_33828;
  wire net_33830;
  wire net_33831;
  wire net_33835;
  wire net_33840;
  wire net_33841;
  wire net_33842;
  wire net_33843;
  wire net_33847;
  wire net_33848;
  wire net_33849;
  wire net_33852;
  wire net_33853;
  wire net_33854;
  wire net_33855;
  wire net_33858;
  wire net_33859;
  wire net_33860;
  wire net_33861;
  wire net_33864;
  wire net_33865;
  wire net_33866;
  wire net_33867;
  wire net_33868;
  wire net_33869;
  wire net_33871;
  wire net_33872;
  wire net_33873;
  wire net_33874;
  wire net_33875;
  wire net_33876;
  wire net_33877;
  wire net_33878;
  wire net_33899;
  wire net_33912;
  wire net_33914;
  wire net_33916;
  wire net_33926;
  wire net_33929;
  wire net_33932;
  wire net_33938;
  wire net_33941;
  wire net_33952;
  wire net_33954;
  wire net_33969;
  wire net_33970;
  wire net_33971;
  wire net_33972;
  wire net_33975;
  wire net_33976;
  wire net_33977;
  wire net_33978;
  wire net_33981;
  wire net_33982;
  wire net_33983;
  wire net_33984;
  wire net_33987;
  wire net_33988;
  wire net_33991;
  wire net_33992;
  wire net_33994;
  wire net_33995;
  wire net_33999;
  wire net_34028;
  wire net_34120;
  wire net_34133;
  wire net_34250;
  wire net_34488;
  wire net_34489;
  wire net_34490;
  wire net_34491;
  wire net_34492;
  wire net_34493;
  wire net_34733;
  wire net_34734;
  wire net_34736;
  wire net_34738;
  wire net_34739;
  wire net_34759;
  wire net_34775;
  wire net_34777;
  wire net_34778;
  wire net_34779;
  wire net_34786;
  wire net_34799;
  wire net_34800;
  wire net_34801;
  wire net_34807;
  wire net_34811;
  wire net_34813;
  wire net_34817;
  wire net_34820;
  wire net_34821;
  wire net_34823;
  wire net_34825;
  wire net_34827;
  wire net_34829;
  wire net_34831;
  wire net_34833;
  wire net_34838;
  wire net_34839;
  wire net_34842;
  wire net_34843;
  wire net_34844;
  wire net_34845;
  wire net_34849;
  wire net_34850;
  wire net_34851;
  wire net_34853;
  wire net_34854;
  wire net_34860;
  wire net_34868;
  wire net_34898;
  wire net_34901;
  wire net_34925;
  wire net_34961;
  wire net_34975;
  wire net_34976;
  wire net_34977;
  wire net_34979;
  wire net_35020;
  wire net_35023;
  wire net_35045;
  wire net_35058;
  wire net_35060;
  wire net_35099;
  wire net_35100;
  wire net_35117;
  wire net_35651;
  wire net_35699;
  wire net_35714;
  wire net_35717;
  wire net_35721;
  wire net_35732;
  wire net_35734;
  wire net_35747;
  wire net_35851;
  wire net_35853;
  wire net_35855;
  wire net_35861;
  wire net_35974;
  wire net_35976;
  wire net_35980;
  wire net_36376;
  wire net_36393;
  wire net_36401;
  wire net_36435;
  wire net_36436;
  wire net_36452;
  wire net_36453;
  wire net_36497;
  wire net_36508;
  wire net_36517;
  wire net_36564;
  wire net_36574;
  wire net_36575;
  wire net_36576;
  wire net_36605;
  wire net_36621;
  wire net_36622;
  wire net_36624;
  wire net_36628;
  wire net_36630;
  wire net_36633;
  wire net_36636;
  wire net_36647;
  wire net_36652;
  wire net_36656;
  wire net_36658;
  wire net_36662;
  wire net_36665;
  wire net_36666;
  wire net_36668;
  wire net_36671;
  wire net_36672;
  wire net_36674;
  wire net_36676;
  wire net_36678;
  wire net_36682;
  wire net_36684;
  wire net_36687;
  wire net_36688;
  wire net_36689;
  wire net_36693;
  wire net_36694;
  wire net_36695;
  wire net_36696;
  wire net_36698;
  wire net_36699;
  wire net_36824;
  wire net_36828;
  wire net_36830;
  wire net_36947;
  wire net_36948;
  wire net_36951;
  wire net_36952;
  wire net_37069;
  wire net_37072;
  wire net_37074;
  wire net_37101;
  wire net_37192;
  wire net_37194;
  wire net_37197;
  wire net_37199;
  wire net_37347;
  wire net_37363;
  wire net_37366;
  wire net_37367;
  wire net_37368;
  wire net_37376;
  wire net_37382;
  wire net_37545;
  wire net_37546;
  wire net_37547;
  wire net_37548;
  wire net_37549;
  wire net_37550;
  wire net_37621;
  wire net_37622;
  wire net_37623;
  wire net_37624;
  wire net_37627;
  wire net_37631;
  wire net_37632;
  wire net_37633;
  wire net_37635;
  wire net_37637;
  wire net_37638;
  wire net_37639;
  wire net_37640;
  wire net_37642;
  wire net_37643;
  wire net_37646;
  wire net_37647;
  wire net_37648;
  wire net_37649;
  wire net_37650;
  wire net_37651;
  wire net_37653;
  wire net_37654;
  wire net_37655;
  wire net_37656;
  wire net_37659;
  wire net_37661;
  wire net_37662;
  wire net_37665;
  wire net_37666;
  wire net_37667;
  wire net_37668;
  wire net_37673;
  wire net_37674;
  wire net_37677;
  wire net_37678;
  wire net_37679;
  wire net_37680;
  wire net_37684;
  wire net_37689;
  wire net_37690;
  wire net_37691;
  wire net_37692;
  wire net_37696;
  wire net_37698;
  wire net_37699;
  wire net_37700;
  wire net_37704;
  wire net_37705;
  wire net_37706;
  wire net_37708;
  wire net_37709;
  wire net_37748;
  wire net_37749;
  wire net_37752;
  wire net_37754;
  wire net_37755;
  wire net_37756;
  wire net_37757;
  wire net_37759;
  wire net_37760;
  wire net_37763;
  wire net_37764;
  wire net_37766;
  wire net_37768;
  wire net_37769;
  wire net_37770;
  wire net_37776;
  wire net_37777;
  wire net_37778;
  wire net_37779;
  wire net_37783;
  wire net_37784;
  wire net_37785;
  wire net_37788;
  wire net_37789;
  wire net_37790;
  wire net_37791;
  wire net_37794;
  wire net_37795;
  wire net_37796;
  wire net_37797;
  wire net_37800;
  wire net_37801;
  wire net_37802;
  wire net_37803;
  wire net_37806;
  wire net_37807;
  wire net_37808;
  wire net_37809;
  wire net_37812;
  wire net_37813;
  wire net_37814;
  wire net_37815;
  wire net_37818;
  wire net_37819;
  wire net_37820;
  wire net_37821;
  wire net_37822;
  wire net_37823;
  wire net_37860;
  wire net_37866;
  wire net_37869;
  wire net_37877;
  wire net_37883;
  wire net_37895;
  wire net_37899;
  wire net_37901;
  wire net_37905;
  wire net_37929;
  wire net_37930;
  wire net_37931;
  wire net_37945;
  wire net_37946;
  wire net_37983;
  wire net_38000;
  wire net_38014;
  wire net_38041;
  wire net_38068;
  wire net_38069;
  wire net_38199;
  wire net_38227;
  wire net_38229;
  wire net_38317;
  wire net_38318;
  wire net_38319;
  wire net_38320;
  wire net_38321;
  wire net_38323;
  wire net_38324;
  wire net_38364;
  wire net_38367;
  wire net_38373;
  wire net_38376;
  wire net_38380;
  wire net_38382;
  wire net_38383;
  wire net_38386;
  wire net_38393;
  wire net_38396;
  wire net_38398;
  wire net_38402;
  wire net_38405;
  wire net_38406;
  wire net_38408;
  wire net_38411;
  wire net_38412;
  wire net_38414;
  wire net_38417;
  wire net_38418;
  wire net_38420;
  wire net_38423;
  wire net_38424;
  wire net_38426;
  wire net_38429;
  wire net_38430;
  wire net_38434;
  wire net_38436;
  wire net_38463;
  wire net_38565;
  wire net_38577;
  wire net_38589;
  wire net_38610;
  wire net_38622;
  wire net_38627;
  wire net_38630;
  wire net_38632;
  wire net_38635;
  wire net_38643;
  wire net_38644;
  wire net_38645;
  wire net_38646;
  wire net_38649;
  wire net_38661;
  wire net_38673;
  wire net_38674;
  wire net_38675;
  wire net_38676;
  wire net_38681;
  wire net_38683;
  wire net_38684;
  wire net_38686;
  wire net_38687;
  wire net_38688;
  wire net_38690;
  wire net_38698;
  wire net_38702;
  wire net_38715;
  wire net_38745;
  wire net_38793;
  wire net_38806;
  wire net_38807;
  wire net_38810;
  wire net_38811;
  wire net_38812;
  wire net_38813;
  wire net_38814;
  wire net_38815;
  wire net_38816;
  wire net_38823;
  wire net_38843;
  wire net_38864;
  wire net_38868;
  wire net_38891;
  wire net_38929;
  wire net_38930;
  wire net_38932;
  wire net_38933;
  wire net_38934;
  wire net_38935;
  wire net_38936;
  wire net_38937;
  wire net_38938;
  wire net_38939;
  wire net_38945;
  wire net_38957;
  wire net_38965;
  wire net_39055;
  wire net_39056;
  wire net_39057;
  wire net_39058;
  wire net_39059;
  wire net_39060;
  wire net_39061;
  wire net_39062;
  wire net_39067;
  wire net_39077;
  wire net_39178;
  wire net_39180;
  wire net_39182;
  wire net_39207;
  wire net_39209;
  wire net_39211;
  wire net_39213;
  wire net_39325;
  wire net_39326;
  wire net_39327;
  wire net_39328;
  wire net_39330;
  wire net_39332;
  wire net_39334;
  wire net_39335;
  wire net_39336;
  wire net_39426;
  wire net_39427;
  wire net_39428;
  wire net_39429;
  wire net_39430;
  wire net_39431;
  wire net_39448;
  wire net_39455;
  wire net_39547;
  wire net_39548;
  wire net_39549;
  wire net_39550;
  wire net_39551;
  wire net_39552;
  wire net_39553;
  wire net_39554;
  wire net_39564;
  wire net_39570;
  wire net_39577;
  wire net_39579;
  wire net_39609;
  wire net_39610;
  wire net_39629;
  wire net_39654;
  wire net_39667;
  wire net_39668;
  wire net_39670;
  wire net_39671;
  wire net_39672;
  wire net_39673;
  wire net_39674;
  wire net_39675;
  wire net_39676;
  wire net_39677;
  wire net_39685;
  wire net_39686;
  wire net_39687;
  wire net_39689;
  wire net_39691;
  wire net_39793;
  wire net_39794;
  wire net_39795;
  wire net_39796;
  wire net_39806;
  wire net_39810;
  wire net_39812;
  wire net_39816;
  wire net_39931;
  wire net_40533;
  wire net_40538;
  wire net_40656;
  wire net_40657;
  wire net_40658;
  wire net_40659;
  wire net_40660;
  wire net_40661;
  wire net_40696;
  wire net_40706;
  wire net_40715;
  wire net_40718;
  wire net_40719;
  wire net_40721;
  wire net_40734;
  wire net_40736;
  wire net_40760;
  wire net_40761;
  wire net_40770;
  wire net_40771;
  wire net_40774;
  wire net_40775;
  wire net_40779;
  wire net_40780;
  wire net_40782;
  wire net_40784;
  wire net_40801;
  wire net_40804;
  wire net_40818;
  wire net_40820;
  wire net_40823;
  wire net_40825;
  wire net_40826;
  wire net_40828;
  wire net_40831;
  wire net_40833;
  wire net_40836;
  wire net_40837;
  wire net_40839;
  wire net_40857;
  wire net_40859;
  wire net_40864;
  wire net_40865;
  wire net_40866;
  wire net_40882;
  wire net_40887;
  wire net_40888;
  wire net_40889;
  wire net_40890;
  wire net_40897;
  wire net_40898;
  wire net_40900;
  wire net_40902;
  wire net_40903;
  wire net_40905;
  wire net_40906;
  wire net_40907;
  wire net_40941;
  wire net_40950;
  wire net_40957;
  wire net_40960;
  wire net_40961;
  wire net_40962;
  wire net_40965;
  wire net_40970;
  wire net_40974;
  wire net_40975;
  wire net_40976;
  wire net_40977;
  wire net_40993;
  wire net_40995;
  wire net_41004;
  wire net_41005;
  wire net_41006;
  wire net_41007;
  wire net_41023;
  wire net_41025;
  wire net_41026;
  wire net_41027;
  wire net_41029;
  wire net_41030;
  wire net_41064;
  wire net_41068;
  wire net_41072;
  wire net_41077;
  wire net_41082;
  wire net_41083;
  wire net_41084;
  wire net_41094;
  wire net_41097;
  wire net_41098;
  wire net_41099;
  wire net_41100;
  wire net_41109;
  wire net_41110;
  wire net_41111;
  wire net_41112;
  wire net_41127;
  wire net_41139;
  wire net_41140;
  wire net_41142;
  wire net_41143;
  wire net_41144;
  wire net_41156;
  wire net_41453;
  wire net_41454;
  wire net_41455;
  wire net_41457;
  wire net_41458;
  wire net_41462;
  wire net_41463;
  wire net_41465;
  wire net_41471;
  wire net_41477;
  wire net_41485;
  wire net_41489;
  wire net_41491;
  wire net_41495;
  wire net_41497;
  wire net_41499;
  wire net_41501;
  wire net_41504;
  wire net_41505;
  wire net_41507;
  wire net_41509;
  wire net_41511;
  wire net_41515;
  wire net_41517;
  wire net_41520;
  wire net_41522;
  wire net_41526;
  wire net_41529;
  wire net_41530;
  wire net_41531;
  wire net_41576;
  wire net_41585;
  wire net_41587;
  wire net_41588;
  wire net_41594;
  wire net_41600;
  wire net_41601;
  wire net_41605;
  wire net_41619;
  wire net_41621;
  wire net_41626;
  wire net_41628;
  wire net_41631;
  wire net_41633;
  wire net_41643;
  wire net_41644;
  wire net_41645;
  wire net_41651;
  wire net_41652;
  wire net_41653;
  wire net_41654;
  wire net_41813;
  wire net_42025;
  wire net_42027;
  wire net_42032;
  wire net_42051;
  wire net_42071;
  wire net_42082;
  wire net_42129;
  wire net_42132;
  wire net_42150;
  wire net_42151;
  wire net_42152;
  wire net_42153;
  wire net_42154;
  wire net_42155;
  wire net_42162;
  wire net_42182;
  wire net_42192;
  wire net_42194;
  wire net_42195;
  wire net_42196;
  wire net_42197;
  wire net_42200;
  wire net_42203;
  wire net_42205;
  wire net_42209;
  wire net_42210;
  wire net_42211;
  wire net_42212;
  wire net_42216;
  wire net_42220;
  wire net_42222;
  wire net_42223;
  wire net_42224;
  wire net_42225;
  wire net_42228;
  wire net_42229;
  wire net_42230;
  wire net_42231;
  wire net_42237;
  wire net_42240;
  wire net_42241;
  wire net_42242;
  wire net_42243;
  wire net_42246;
  wire net_42258;
  wire net_42264;
  wire net_42265;
  wire net_42266;
  wire net_42267;
  wire net_42268;
  wire net_42269;
  wire net_42271;
  wire net_42272;
  wire net_42274;
  wire net_42275;
  wire net_42276;
  wire net_42277;
  wire net_42278;
  wire net_42295;
  wire net_42394;
  wire net_42397;
  wire net_42398;
  wire net_42399;
  wire net_42400;
  wire net_42401;
  wire net_42409;
  wire net_42413;
  wire net_42419;
  wire net_42436;
  wire net_42441;
  wire net_42481;
  wire net_42482;
  wire net_42519;
  wire net_42524;
  wire net_42530;
  wire net_42534;
  wire net_42535;
  wire net_42545;
  wire net_42549;
  wire net_42560;
  wire net_42563;
  wire net_42576;
  wire net_42578;
  wire net_42581;
  wire net_42586;
  wire net_42587;
  wire net_42593;
  wire net_42597;
  wire net_42603;
  wire net_42605;
  wire net_42606;
  wire net_42618;
  wire net_42637;
  wire net_42638;
  wire net_42641;
  wire net_42642;
  wire net_42643;
  wire net_42644;
  wire net_42646;
  wire net_42647;
  wire net_42665;
  wire net_42674;
  wire net_42681;
  wire net_42682;
  wire net_42684;
  wire net_42685;
  wire net_42686;
  wire net_42687;
  wire net_42689;
  wire net_42690;
  wire net_42692;
  wire net_42693;
  wire net_42696;
  wire net_42698;
  wire net_42699;
  wire net_42700;
  wire net_42702;
  wire net_42703;
  wire net_42708;
  wire net_42713;
  wire net_42715;
  wire net_42716;
  wire net_42719;
  wire net_42721;
  wire net_42722;
  wire net_42723;
  wire net_42725;
  wire net_42727;
  wire net_42728;
  wire net_42729;
  wire net_42731;
  wire net_42733;
  wire net_42734;
  wire net_42735;
  wire net_42737;
  wire net_42739;
  wire net_42740;
  wire net_42741;
  wire net_42743;
  wire net_42745;
  wire net_42746;
  wire net_42747;
  wire net_42749;
  wire net_42751;
  wire net_42752;
  wire net_42753;
  wire net_42755;
  wire net_42757;
  wire net_42758;
  wire net_42759;
  wire net_42760;
  wire net_42761;
  wire net_42763;
  wire net_42764;
  wire net_42765;
  wire net_42766;
  wire net_42767;
  wire net_42768;
  wire net_42769;
  wire net_42770;
  wire net_42778;
  wire net_42780;
  wire net_42781;
  wire net_42783;
  wire net_42785;
  wire net_42786;
  wire net_42794;
  wire net_42799;
  wire net_42804;
  wire net_42805;
  wire net_42807;
  wire net_42808;
  wire net_42809;
  wire net_42810;
  wire net_42811;
  wire net_42812;
  wire net_42813;
  wire net_42815;
  wire net_42817;
  wire net_42822;
  wire net_42823;
  wire net_42828;
  wire net_42831;
  wire net_42832;
  wire net_42835;
  wire net_42836;
  wire net_42838;
  wire net_42839;
  wire net_42840;
  wire net_42842;
  wire net_42844;
  wire net_42845;
  wire net_42846;
  wire net_42848;
  wire net_42850;
  wire net_42851;
  wire net_42852;
  wire net_42854;
  wire net_42856;
  wire net_42857;
  wire net_42858;
  wire net_42860;
  wire net_42862;
  wire net_42863;
  wire net_42864;
  wire net_42866;
  wire net_42868;
  wire net_42869;
  wire net_42870;
  wire net_42872;
  wire net_42874;
  wire net_42875;
  wire net_42876;
  wire net_42880;
  wire net_42881;
  wire net_42882;
  wire net_42883;
  wire net_42884;
  wire net_42886;
  wire net_42887;
  wire net_42888;
  wire net_42889;
  wire net_42890;
  wire net_42891;
  wire net_42892;
  wire net_42893;
  wire net_42895;
  wire net_42898;
  wire net_42899;
  wire net_42906;
  wire net_42909;
  wire net_42927;
  wire net_42936;
  wire net_42938;
  wire net_42941;
  wire net_42942;
  wire net_42945;
  wire net_42947;
  wire net_42958;
  wire net_42962;
  wire net_42969;
  wire net_42974;
  wire net_42981;
  wire net_42984;
  wire net_42992;
  wire net_42998;
  wire net_43003;
  wire net_43006;
  wire net_43007;
  wire net_43011;
  wire net_43012;
  wire net_43013;
  wire net_43015;
  wire net_43026;
  wire net_43027;
  wire net_43037;
  wire net_43041;
  wire net_43043;
  wire net_43052;
  wire net_43056;
  wire net_43074;
  wire net_43085;
  wire net_43096;
  wire net_43109;
  wire net_43129;
  wire net_43130;
  wire net_43137;
  wire net_43150;
  wire net_43152;
  wire net_43156;
  wire net_43157;
  wire net_43158;
  wire net_43159;
  wire net_43160;
  wire net_43162;
  wire net_43164;
  wire net_43166;
  wire net_43256;
  wire net_43279;
  wire net_43280;
  wire net_43281;
  wire net_43282;
  wire net_43283;
  wire net_43285;
  wire net_43286;
  wire net_43290;
  wire net_43300;
  wire net_43302;
  wire net_43309;
  wire net_43311;
  wire net_43315;
  wire net_43321;
  wire net_43322;
  wire net_43325;
  wire net_43331;
  wire net_43334;
  wire net_43336;
  wire net_43340;
  wire net_43342;
  wire net_43344;
  wire net_43346;
  wire net_43349;
  wire net_43350;
  wire net_43352;
  wire net_43355;
  wire net_43356;
  wire net_43358;
  wire net_43360;
  wire net_43362;
  wire net_43364;
  wire net_43367;
  wire net_43368;
  wire net_43370;
  wire net_43372;
  wire net_43374;
  wire net_43376;
  wire net_43379;
  wire net_43380;
  wire net_43381;
  wire net_43382;
  wire net_43383;
  wire net_43398;
  wire net_43399;
  wire net_43400;
  wire net_43403;
  wire net_43405;
  wire net_43407;
  wire net_43408;
  wire net_43411;
  wire net_43413;
  wire net_43414;
  wire net_43424;
  wire net_43430;
  wire net_43436;
  wire net_43437;
  wire net_43441;
  wire net_43443;
  wire net_43447;
  wire net_43450;
  wire net_43451;
  wire net_43453;
  wire net_43455;
  wire net_43457;
  wire net_43460;
  wire net_43461;
  wire net_43463;
  wire net_43466;
  wire net_43467;
  wire net_43469;
  wire net_43471;
  wire net_43473;
  wire net_43475;
  wire net_43477;
  wire net_43479;
  wire net_43481;
  wire net_43484;
  wire net_43485;
  wire net_43487;
  wire net_43490;
  wire net_43491;
  wire net_43493;
  wire net_43495;
  wire net_43497;
  wire net_43499;
  wire net_43503;
  wire net_43504;
  wire net_43507;
  wire net_43519;
  wire net_43523;
  wire net_43526;
  wire net_43528;
  wire net_43532;
  wire net_43534;
  wire net_43537;
  wire net_43544;
  wire net_43548;
  wire net_43549;
  wire net_43550;
  wire net_43551;
  wire net_43554;
  wire net_43569;
  wire net_43571;
  wire net_43574;
  wire net_43576;
  wire net_43578;
  wire net_43580;
  wire net_43582;
  wire net_43584;
  wire net_43586;
  wire net_43589;
  wire net_43590;
  wire net_43592;
  wire net_43594;
  wire net_43596;
  wire net_43598;
  wire net_43600;
  wire net_43602;
  wire net_43604;
  wire net_43606;
  wire net_43608;
  wire net_43610;
  wire net_43613;
  wire net_43614;
  wire net_43616;
  wire net_43619;
  wire net_43620;
  wire net_43622;
  wire net_43625;
  wire net_43626;
  wire net_43630;
  wire net_43636;
  wire net_43638;
  wire net_43640;
  wire net_43642;
  wire net_43644;
  wire net_43646;
  wire net_43660;
  wire net_43666;
  wire net_43668;
  wire net_43673;
  wire net_43691;
  wire net_43697;
  wire net_43699;
  wire net_43701;
  wire net_43703;
  wire net_43706;
  wire net_43707;
  wire net_43709;
  wire net_43711;
  wire net_43713;
  wire net_43718;
  wire net_43719;
  wire net_43745;
  wire net_43759;
  wire net_43760;
  wire net_43763;
  wire net_43765;
  wire net_43767;
  wire net_43892;
  wire net_43999;
  wire net_44138;
  wire net_44148;
  wire net_44250;
  wire net_44413;
  wire net_44430;
  wire net_44434;
  wire net_44448;
  wire net_44451;
  wire net_44478;
  wire net_44482;
  wire net_44483;
  wire net_44520;
  wire net_44529;
  wire net_44531;
  wire net_44532;
  wire net_44533;
  wire net_44537;
  wire net_44539;
  wire net_44541;
  wire net_44549;
  wire net_44553;
  wire net_44554;
  wire net_44561;
  wire net_44564;
  wire net_44567;
  wire net_44570;
  wire net_44572;
  wire net_44574;
  wire net_44576;
  wire net_44579;
  wire net_44580;
  wire net_44582;
  wire net_44584;
  wire net_44586;
  wire net_44590;
  wire net_44592;
  wire net_44595;
  wire net_44596;
  wire net_44601;
  wire net_44604;
  wire net_44605;
  wire net_44606;
  wire net_44653;
  wire net_44655;
  wire net_44656;
  wire net_44660;
  wire net_44663;
  wire net_44664;
  wire net_44670;
  wire net_44675;
  wire net_44676;
  wire net_44680;
  wire net_44694;
  wire net_44695;
  wire net_44696;
  wire net_44697;
  wire net_44701;
  wire net_44702;
  wire net_44703;
  wire net_44712;
  wire net_44713;
  wire net_44714;
  wire net_44715;
  wire net_44726;
  wire net_44727;
  wire net_44728;
  wire net_44729;
  wire net_44736;
  wire net_44773;
  wire net_44774;
  wire net_44783;
  wire net_44784;
  wire net_44788;
  wire net_44793;
  wire net_44803;
  wire net_44805;
  wire net_44806;
  wire net_44807;
  wire net_44808;
  wire net_44817;
  wire net_44818;
  wire net_44823;
  wire net_44824;
  wire net_44825;
  wire net_44826;
  wire net_44835;
  wire net_44836;
  wire net_44837;
  wire net_44838;
  wire net_44841;
  wire net_44842;
  wire net_44843;
  wire net_44844;
  wire net_44847;
  wire net_44848;
  wire net_44849;
  wire net_44850;
  wire net_44851;
  wire net_44852;
  wire net_44855;
  wire net_44857;
  wire net_44895;
  wire net_44897;
  wire net_44899;
  wire net_44900;
  wire net_44903;
  wire net_44905;
  wire net_44907;
  wire net_44908;
  wire net_44911;
  wire net_44913;
  wire net_44917;
  wire net_44922;
  wire net_44923;
  wire net_44925;
  wire net_44926;
  wire net_44929;
  wire net_44930;
  wire net_44940;
  wire net_44941;
  wire net_44942;
  wire net_44943;
  wire net_44946;
  wire net_44947;
  wire net_44948;
  wire net_44949;
  wire net_44952;
  wire net_44953;
  wire net_44954;
  wire net_44955;
  wire net_44964;
  wire net_44965;
  wire net_44966;
  wire net_44967;
  wire net_44970;
  wire net_44971;
  wire net_44972;
  wire net_44973;
  wire net_44974;
  wire net_44975;
  wire net_45762;
  wire net_45907;
  wire net_45908;
  wire net_45911;
  wire net_45912;
  wire net_45921;
  wire net_45923;
  wire net_45924;
  wire net_45930;
  wire net_45931;
  wire net_45932;
  wire net_45933;
  wire net_45943;
  wire net_45945;
  wire net_45972;
  wire net_45974;
  wire net_45976;
  wire net_45977;
  wire net_45980;
  wire net_45984;
  wire net_45985;
  wire net_46011;
  wire net_46020;
  wire net_46021;
  wire net_46022;
  wire net_46023;
  wire net_46024;
  wire net_46028;
  wire net_46030;
  wire net_46034;
  wire net_46035;
  wire net_46037;
  wire net_46054;
  wire net_46058;
  wire net_46060;
  wire net_46061;
  wire net_46064;
  wire net_46066;
  wire net_46067;
  wire net_46068;
  wire net_46070;
  wire net_46072;
  wire net_46073;
  wire net_46074;
  wire net_46076;
  wire net_46078;
  wire net_46079;
  wire net_46080;
  wire net_46082;
  wire net_46084;
  wire net_46085;
  wire net_46086;
  wire net_46088;
  wire net_46090;
  wire net_46091;
  wire net_46092;
  wire net_46095;
  wire net_46097;
  wire net_46098;
  wire net_46127;
  wire net_46145;
  wire net_46146;
  wire net_46147;
  wire net_46148;
  wire net_46149;
  wire net_46150;
  wire net_46154;
  wire net_46155;
  wire net_46156;
  wire net_46157;
  wire net_46158;
  wire net_46165;
  wire net_46167;
  wire net_46179;
  wire net_46183;
  wire net_46197;
  wire net_46200;
  wire net_46201;
  wire net_46202;
  wire net_46203;
  wire net_46206;
  wire net_46207;
  wire net_46208;
  wire net_46209;
  wire net_46212;
  wire net_46213;
  wire net_46214;
  wire net_46215;
  wire net_46218;
  wire net_46219;
  wire net_46220;
  wire net_46221;
  wire net_46222;
  wire net_46223;
  wire net_46249;
  wire net_46253;
  wire net_46255;
  wire net_46257;
  wire net_46268;
  wire net_46269;
  wire net_46271;
  wire net_46273;
  wire net_46276;
  wire net_46277;
  wire net_46279;
  wire net_46286;
  wire net_46292;
  wire net_46294;
  wire net_46297;
  wire net_46299;
  wire net_46300;
  wire net_46301;
  wire net_46302;
  wire net_46317;
  wire net_46319;
  wire net_46324;
  wire net_46329;
  wire net_46331;
  wire net_46336;
  wire net_46337;
  wire net_46338;
  wire net_46341;
  wire net_46342;
  wire net_46345;
  wire net_46346;
  wire net_46347;
  wire net_46348;
  wire net_46349;
  wire net_46350;
  wire net_46351;
  wire net_46353;
  wire net_46354;
  wire net_46363;
  wire net_46370;
  wire net_46375;
  wire net_46377;
  wire net_46383;
  wire net_46407;
  wire net_46419;
  wire net_46436;
  wire net_46464;
  wire net_46468;
  wire net_46469;
  wire net_46472;
  wire net_46473;
  wire net_46474;
  wire net_46475;
  wire net_46476;
  wire net_46477;
  wire net_46478;
  wire net_46504;
  wire net_46513;
  wire net_46514;
  wire net_46517;
  wire net_46519;
  wire net_46525;
  wire net_46529;
  wire net_46532;
  wire net_46533;
  wire net_46534;
  wire net_46535;
  wire net_46537;
  wire net_46551;
  wire net_46552;
  wire net_46553;
  wire net_46554;
  wire net_46557;
  wire net_46563;
  wire net_46564;
  wire net_46565;
  wire net_46566;
  wire net_46569;
  wire net_46570;
  wire net_46571;
  wire net_46572;
  wire net_46581;
  wire net_46588;
  wire net_46591;
  wire net_46592;
  wire net_46594;
  wire net_46595;
  wire net_46596;
  wire net_46597;
  wire net_46598;
  wire net_46599;
  wire net_46600;
  wire net_46601;
  wire net_46610;
  wire net_46612;
  wire net_46613;
  wire net_46614;
  wire net_46615;
  wire net_46616;
  wire net_46625;
  wire net_46639;
  wire net_46640;
  wire net_46641;
  wire net_46642;
  wire net_46644;
  wire net_46645;
  wire net_46646;
  wire net_46647;
  wire net_46648;
  wire net_46650;
  wire net_46652;
  wire net_46653;
  wire net_46656;
  wire net_46658;
  wire net_46663;
  wire net_46665;
  wire net_46668;
  wire net_46669;
  wire net_46670;
  wire net_46671;
  wire net_46674;
  wire net_46675;
  wire net_46676;
  wire net_46677;
  wire net_46680;
  wire net_46681;
  wire net_46682;
  wire net_46683;
  wire net_46688;
  wire net_46692;
  wire net_46693;
  wire net_46694;
  wire net_46695;
  wire net_46698;
  wire net_46699;
  wire net_46700;
  wire net_46701;
  wire net_46704;
  wire net_46705;
  wire net_46706;
  wire net_46707;
  wire net_46712;
  wire net_46717;
  wire net_46718;
  wire net_46719;
  wire net_46720;
  wire net_46721;
  wire net_46722;
  wire net_46724;
  wire net_46733;
  wire net_46735;
  wire net_46737;
  wire net_46743;
  wire net_46751;
  wire net_46758;
  wire net_46760;
  wire net_46762;
  wire net_46764;
  wire net_46765;
  wire net_46768;
  wire net_46769;
  wire net_46773;
  wire net_46774;
  wire net_46776;
  wire net_46780;
  wire net_46784;
  wire net_46794;
  wire net_46798;
  wire net_46800;
  wire net_46805;
  wire net_46812;
  wire net_46815;
  wire net_46821;
  wire net_46822;
  wire net_46823;
  wire net_46824;
  wire net_46829;
  wire net_46833;
  wire net_46834;
  wire net_46835;
  wire net_46836;
  wire net_46837;
  wire net_46838;
  wire net_46840;
  wire net_46841;
  wire net_46842;
  wire net_46843;
  wire net_46844;
  wire net_46845;
  wire net_46847;
  wire net_46856;
  wire net_46857;
  wire net_46884;
  wire net_46892;
  wire net_46894;
  wire net_46898;
  wire net_46905;
  wire net_46927;
  wire net_46932;
  wire net_46940;
  wire net_46951;
  wire net_46960;
  wire net_46961;
  wire net_46964;
  wire net_46965;
  wire net_46967;
  wire net_46968;
  wire net_46969;
  wire net_46979;
  wire net_47006;
  wire net_47009;
  wire net_47069;
  wire net_47083;
  wire net_47084;
  wire net_47086;
  wire net_47087;
  wire net_47089;
  wire net_47091;
  wire net_47092;
  wire net_47100;
  wire net_47102;
  wire net_47117;
  wire net_47120;
  wire net_47128;
  wire net_47148;
  wire net_47166;
  wire net_47168;
  wire net_47207;
  wire net_47209;
  wire net_47211;
  wire net_47214;
  wire net_47216;
  wire net_47225;
  wire net_47252;
  wire net_47258;
  wire net_47268;
  wire net_47269;
  wire net_47271;
  wire net_47272;
  wire net_47274;
  wire net_47275;
  wire net_47276;
  wire net_47279;
  wire net_47289;
  wire net_47290;
  wire net_47291;
  wire net_47292;
  wire net_47295;
  wire net_47296;
  wire net_47297;
  wire net_47298;
  wire net_47304;
  wire net_47308;
  wire net_47314;
  wire net_47329;
  wire net_47330;
  wire net_47334;
  wire net_47335;
  wire net_47336;
  wire net_47338;
  wire net_47339;
  wire net_47348;
  wire net_47350;
  wire net_47351;
  wire net_47357;
  wire net_47361;
  wire net_47365;
  wire net_47374;
  wire net_47377;
  wire net_47382;
  wire net_47385;
  wire net_47391;
  wire net_47397;
  wire net_47403;
  wire net_47418;
  wire net_47419;
  wire net_47420;
  wire net_47421;
  wire net_47424;
  wire net_47445;
  wire net_47452;
  wire net_47453;
  wire net_47456;
  wire net_47475;
  wire net_47483;
  wire net_47498;
  wire net_47505;
  wire net_47516;
  wire net_47538;
  wire net_47543;
  wire net_47565;
  wire net_47575;
  wire net_47576;
  wire net_47578;
  wire net_47580;
  wire net_47582;
  wire net_47584;
  wire net_47585;
  wire net_47596;
  wire net_47603;
  wire net_47718;
  wire net_47720;
  wire net_47724;
  wire net_47726;
  wire net_47824;
  wire net_47883;
  wire net_47892;
  wire net_47936;
  wire net_47944;
  wire net_47945;
  wire net_48318;
  wire net_48319;
  wire net_48320;
  wire net_48321;
  wire net_48322;
  wire net_48323;
  wire net_48440;
  wire net_48441;
  wire net_48452;
  wire net_48456;
  wire net_48583;
  wire net_48606;
  wire net_48616;
  wire net_48668;
  wire net_48669;
  wire net_48691;
  wire net_48737;
  wire net_48738;
  wire net_48742;
  wire net_48747;
  wire net_48765;
  wire net_48766;
  wire net_48767;
  wire net_48768;
  wire net_48777;
  wire net_48778;
  wire net_48779;
  wire net_48780;
  wire net_48810;
  wire net_48817;
  wire net_48824;
  wire net_49196;
  wire net_49202;
  wire net_49320;
  wire net_49321;
  wire net_49322;
  wire net_49323;
  wire net_49324;
  wire net_49325;
  wire net_49700;
  wire net_49812;
  wire net_49813;
  wire net_49814;
  wire net_49815;
  wire net_49816;
  wire net_49817;
  wire net_49862;
  wire net_49866;
  wire net_49872;
  wire net_49875;
  wire net_49876;
  wire net_49880;
  wire net_49892;
  wire net_49915;
  wire net_49920;
  wire net_49922;
  wire net_49923;
  wire net_49930;
  wire net_49931;
  wire net_49933;
  wire net_49934;
  wire net_49935;
  wire net_49938;
  wire net_49939;
  wire net_49946;
  wire net_49949;
  wire net_50091;
  wire net_50180;
  wire net_50185;
  wire net_50220;
  wire net_50223;
  wire net_50226;
  wire net_50227;
  wire net_50229;
  wire net_50230;
  wire net_50234;
  wire net_50239;
  wire net_50240;
  wire net_50247;
  wire net_50253;
  wire net_50259;
  wire net_50260;
  wire net_50261;
  wire net_50262;
  wire net_50265;
  wire net_50271;
  wire net_50272;
  wire net_50273;
  wire net_50274;
  wire net_50284;
  wire net_50292;
  wire net_50299;
  wire net_50300;
  wire net_50302;
  wire net_50303;
  wire net_50304;
  wire net_50305;
  wire net_50306;
  wire net_50307;
  wire net_50308;
  wire net_50309;
  wire net_50313;
  wire net_50318;
  wire net_50343;
  wire net_50344;
  wire net_50345;
  wire net_50346;
  wire net_50347;
  wire net_50348;
  wire net_50349;
  wire net_50351;
  wire net_50353;
  wire net_50354;
  wire net_50355;
  wire net_50356;
  wire net_50359;
  wire net_50360;
  wire net_50361;
  wire net_50370;
  wire net_50371;
  wire net_50375;
  wire net_50377;
  wire net_50378;
  wire net_50381;
  wire net_50383;
  wire net_50384;
  wire net_50385;
  wire net_50387;
  wire net_50389;
  wire net_50390;
  wire net_50391;
  wire net_50393;
  wire net_50395;
  wire net_50396;
  wire net_50397;
  wire net_50399;
  wire net_50401;
  wire net_50402;
  wire net_50403;
  wire net_50405;
  wire net_50407;
  wire net_50408;
  wire net_50409;
  wire net_50411;
  wire net_50413;
  wire net_50414;
  wire net_50415;
  wire net_50417;
  wire net_50419;
  wire net_50420;
  wire net_50421;
  wire net_50422;
  wire net_50423;
  wire net_50425;
  wire net_50426;
  wire net_50427;
  wire net_50428;
  wire net_50429;
  wire net_50430;
  wire net_50431;
  wire net_50432;
  wire net_50443;
  wire net_50451;
  wire net_50461;
  wire net_50466;
  wire net_50467;
  wire net_50468;
  wire net_50469;
  wire net_50471;
  wire net_50474;
  wire net_50475;
  wire net_50477;
  wire net_50478;
  wire net_50479;
  wire net_50481;
  wire net_50483;
  wire net_50484;
  wire net_50485;
  wire net_50492;
  wire net_50493;
  wire net_50495;
  wire net_50498;
  wire net_50500;
  wire net_50501;
  wire net_50502;
  wire net_50504;
  wire net_50506;
  wire net_50507;
  wire net_50508;
  wire net_50510;
  wire net_50512;
  wire net_50513;
  wire net_50514;
  wire net_50516;
  wire net_50518;
  wire net_50519;
  wire net_50520;
  wire net_50522;
  wire net_50524;
  wire net_50525;
  wire net_50526;
  wire net_50528;
  wire net_50530;
  wire net_50531;
  wire net_50532;
  wire net_50534;
  wire net_50536;
  wire net_50537;
  wire net_50538;
  wire net_50542;
  wire net_50543;
  wire net_50544;
  wire net_50545;
  wire net_50546;
  wire net_50548;
  wire net_50549;
  wire net_50550;
  wire net_50551;
  wire net_50552;
  wire net_50553;
  wire net_50554;
  wire net_50555;
  wire net_50560;
  wire net_50564;
  wire net_50567;
  wire net_50568;
  wire net_50570;
  wire net_50593;
  wire net_50597;
  wire net_50598;
  wire net_50599;
  wire net_50600;
  wire net_50601;
  wire net_50602;
  wire net_50603;
  wire net_50609;
  wire net_50613;
  wire net_50615;
  wire net_50616;
  wire net_50617;
  wire net_50620;
  wire net_50622;
  wire net_50623;
  wire net_50624;
  wire net_50631;
  wire net_50634;
  wire net_50635;
  wire net_50636;
  wire net_50637;
  wire net_50640;
  wire net_50649;
  wire net_50654;
  wire net_50664;
  wire net_50665;
  wire net_50666;
  wire net_50667;
  wire net_50668;
  wire net_50669;
  wire net_50671;
  wire net_50672;
  wire net_50673;
  wire net_50674;
  wire net_50675;
  wire net_50676;
  wire net_50677;
  wire net_50678;
  wire net_50689;
  wire net_50697;
  wire net_50698;
  wire net_50712;
  wire net_50713;
  wire net_50716;
  wire net_50718;
  wire net_50722;
  wire net_50724;
  wire net_50726;
  wire net_50728;
  wire net_50735;
  wire net_50740;
  wire net_50743;
  wire net_50745;
  wire net_50752;
  wire net_50757;
  wire net_50758;
  wire net_50759;
  wire net_50760;
  wire net_50763;
  wire net_50769;
  wire net_50770;
  wire net_50771;
  wire net_50772;
  wire net_50775;
  wire net_50776;
  wire net_50777;
  wire net_50778;
  wire net_50789;
  wire net_50791;
  wire net_50792;
  wire net_50795;
  wire net_50796;
  wire net_50797;
  wire net_50798;
  wire net_50799;
  wire net_50800;
  wire net_50801;
  wire net_50811;
  wire net_50812;
  wire net_50813;
  wire net_50835;
  wire net_50836;
  wire net_50854;
  wire net_50861;
  wire net_50862;
  wire net_50865;
  wire net_50876;
  wire net_50883;
  wire net_50893;
  wire net_50898;
  wire net_50899;
  wire net_50905;
  wire net_50906;
  wire net_50914;
  wire net_50915;
  wire net_50917;
  wire net_50918;
  wire net_50919;
  wire net_50920;
  wire net_50921;
  wire net_50922;
  wire net_50923;
  wire net_50924;
  wire net_50939;
  wire net_50960;
  wire net_50962;
  wire net_50963;
  wire net_50967;
  wire net_50971;
  wire net_50980;
  wire net_50993;
  wire net_50999;
  wire net_51012;
  wire net_51022;
  wire net_51027;
  wire net_51037;
  wire net_51038;
  wire net_51043;
  wire net_51044;
  wire net_51045;
  wire net_51054;
  wire net_51055;
  wire net_51059;
  wire net_51063;
  wire net_51071;
  wire net_51082;
  wire net_51085;
  wire net_51086;
  wire net_51088;
  wire net_51095;
  wire net_51099;
  wire net_51101;
  wire net_51103;
  wire net_51105;
  wire net_51106;
  wire net_51114;
  wire net_51115;
  wire net_51116;
  wire net_51117;
  wire net_51126;
  wire net_51127;
  wire net_51128;
  wire net_51129;
  wire net_51144;
  wire net_51157;
  wire net_51160;
  wire net_51161;
  wire net_51164;
  wire net_51165;
  wire net_51167;
  wire net_51169;
  wire net_51170;
  wire net_51175;
  wire net_51187;
  wire net_51191;
  wire net_51195;
  wire net_51210;
  wire net_51213;
  wire net_51214;
  wire net_51215;
  wire net_51216;
  wire net_51220;
  wire net_51222;
  wire net_51228;
  wire net_51231;
  wire net_51235;
  wire net_51249;
  wire net_51250;
  wire net_51251;
  wire net_51252;
  wire net_51256;
  wire net_51261;
  wire net_51263;
  wire net_51276;
  wire net_51280;
  wire net_51282;
  wire net_51283;
  wire net_51284;
  wire net_51286;
  wire net_51287;
  wire net_51289;
  wire net_51290;
  wire net_51291;
  wire net_51292;
  wire net_51293;
  wire net_51303;
  wire net_51304;
  wire net_51307;
  wire net_51310;
  wire net_51311;
  wire net_51315;
  wire net_51319;
  wire net_51343;
  wire net_51367;
  wire net_51406;
  wire net_51407;
  wire net_51415;
  wire net_51432;
  wire net_51433;
  wire net_51452;
  wire net_51456;
  wire net_51460;
  wire net_51461;
  wire net_51470;
  wire net_51471;
  wire net_51473;
  wire net_51477;
  wire net_51484;
  wire net_51485;
  wire net_51498;
  wire net_51508;
  wire net_51510;
  wire net_51521;
  wire net_51522;
  wire net_51525;
  wire net_51526;
  wire net_51527;
  wire net_51528;
  wire net_51529;
  wire net_51530;
  wire net_51531;
  wire net_51533;
  wire net_51535;
  wire net_51537;
  wire net_51539;
  wire net_51543;
  wire net_51544;
  wire net_51550;
  wire net_51555;
  wire net_51681;
  wire net_51719;
  wire net_51730;
  wire net_51776;
  wire net_51799;
  wire net_52149;
  wire net_52151;
  wire net_52152;
  wire net_52153;
  wire net_52154;
  wire net_52195;
  wire net_52197;
  wire net_52199;
  wire net_52206;
  wire net_52207;
  wire net_52208;
  wire net_52209;
  wire net_52211;
  wire net_52215;
  wire net_52218;
  wire net_52223;
  wire net_52226;
  wire net_52229;
  wire net_52232;
  wire net_52234;
  wire net_52236;
  wire net_52238;
  wire net_52241;
  wire net_52242;
  wire net_52244;
  wire net_52246;
  wire net_52248;
  wire net_52252;
  wire net_52254;
  wire net_52257;
  wire net_52258;
  wire net_52264;
  wire net_52266;
  wire net_52267;
  wire net_52268;
  wire net_52313;
  wire net_52320;
  wire net_52321;
  wire net_52322;
  wire net_52336;
  wire net_52352;
  wire net_52353;
  wire net_52356;
  wire net_52358;
  wire net_52390;
  wire net_52391;
  wire net_52407;
  wire net_52408;
  wire net_52639;
  wire net_52640;
  wire net_52679;
  wire net_52869;
  wire net_52870;
  wire net_52872;
  wire net_52873;
  wire net_52929;
  wire net_53026;
  wire net_53027;
  wire net_53028;
  wire net_53029;
  wire net_53030;
  wire net_53031;
  wire net_53032;
  wire net_53033;
  wire net_53073;
  wire net_53074;
  wire net_53078;
  wire net_53092;
  wire net_53095;
  wire net_53098;
  wire net_53109;
  wire net_53142;
  wire net_53143;
  wire net_53144;
  wire net_53145;
  wire net_53146;
  wire net_53147;
  wire net_53149;
  wire net_53150;
  wire net_53151;
  wire net_53153;
  wire net_53154;
  wire net_53156;
  wire net_53194;
  wire net_53198;
  wire net_53204;
  wire net_53208;
  wire net_53210;
  wire net_53211;
  wire net_53213;
  wire net_53214;
  wire net_53215;
  wire net_53221;
  wire net_53225;
  wire net_53228;
  wire net_53231;
  wire net_53234;
  wire net_53237;
  wire net_53238;
  wire net_53240;
  wire net_53242;
  wire net_53244;
  wire net_53246;
  wire net_53248;
  wire net_53250;
  wire net_53255;
  wire net_53256;
  wire net_53259;
  wire net_53260;
  wire net_53265;
  wire net_53267;
  wire net_53269;
  wire net_53270;
  wire net_53519;
  wire net_53524;
  wire net_53525;
  wire net_53547;
  wire net_53645;
  wire net_53646;
  wire net_53647;
  wire net_53648;
  wire net_53674;
  wire net_53682;
  wire net_53683;
  wire net_53687;
  wire net_53688;
  wire net_53690;
  wire net_53696;
  wire net_53712;
  wire net_53713;
  wire net_53716;
  wire net_53720;
  wire net_53722;
  wire net_53726;
  wire net_53728;
  wire net_53730;
  wire net_53732;
  wire net_53735;
  wire net_53736;
  wire net_53738;
  wire net_53741;
  wire net_53742;
  wire net_53744;
  wire net_53747;
  wire net_53748;
  wire net_53750;
  wire net_53753;
  wire net_53754;
  wire net_53759;
  wire net_53760;
  wire net_53766;
  wire net_53767;
  wire net_53768;
  wire net_53769;
  wire net_53770;
  wire net_53771;
  wire net_53786;
  wire net_53807;
  wire net_53809;
  wire net_53814;
  wire net_53815;
  wire net_53817;
  wire net_53818;
  wire net_53819;
  wire net_53820;
  wire net_53823;
  wire net_53825;
  wire net_53827;
  wire net_53831;
  wire net_53832;
  wire net_53834;
  wire net_53836;
  wire net_53838;
  wire net_53839;
  wire net_53840;
  wire net_53841;
  wire net_53844;
  wire net_53845;
  wire net_53846;
  wire net_53847;
  wire net_53850;
  wire net_53851;
  wire net_53852;
  wire net_53853;
  wire net_53868;
  wire net_53869;
  wire net_53870;
  wire net_53871;
  wire net_53874;
  wire net_53875;
  wire net_53876;
  wire net_53877;
  wire net_53884;
  wire net_53885;
  wire net_53894;
  wire net_54010;
  wire net_54011;
  wire net_54012;
  wire net_54013;
  wire net_54014;
  wire net_54015;
  wire net_54016;
  wire net_54017;
  wire net_54022;
  wire net_54064;
  wire net_54069;
  wire net_54081;
  wire net_54090;
  wire net_54120;
  wire net_54130;
  wire net_54131;
  wire net_54133;
  wire net_54134;
  wire net_54135;
  wire net_54136;
  wire net_54137;
  wire net_54138;
  wire net_54139;
  wire net_54140;
  wire net_54157;
  wire net_54159;
  wire net_54161;
  wire net_54162;
  wire net_54166;
  wire net_54175;
  wire net_54176;
  wire net_54177;
  wire net_54178;
  wire net_54179;
  wire net_54186;
  wire net_54187;
  wire net_54188;
  wire net_54189;
  wire net_54190;
  wire net_54191;
  wire net_54193;
  wire net_54195;
  wire net_54202;
  wire net_54205;
  wire net_54207;
  wire net_54208;
  wire net_54209;
  wire net_54210;
  wire net_54214;
  wire net_54215;
  wire net_54219;
  wire net_54220;
  wire net_54221;
  wire net_54222;
  wire net_54225;
  wire net_54226;
  wire net_54227;
  wire net_54228;
  wire net_54234;
  wire net_54238;
  wire net_54243;
  wire net_54244;
  wire net_54245;
  wire net_54246;
  wire net_54252;
  wire net_54253;
  wire net_54254;
  wire net_54256;
  wire net_54257;
  wire net_54258;
  wire net_54259;
  wire net_54260;
  wire net_54261;
  wire net_54262;
  wire net_54263;
  wire net_54268;
  wire net_54275;
  wire net_54276;
  wire net_54281;
  wire net_54282;
  wire net_54283;
  wire net_54285;
  wire net_54288;
  wire net_54291;
  wire net_54297;
  wire net_54299;
  wire net_54300;
  wire net_54302;
  wire net_54305;
  wire net_54308;
  wire net_54309;
  wire net_54310;
  wire net_54312;
  wire net_54316;
  wire net_54318;
  wire net_54319;
  wire net_54323;
  wire net_54325;
  wire net_54326;
  wire net_54328;
  wire net_54330;
  wire net_54331;
  wire net_54332;
  wire net_54333;
  wire net_54338;
  wire net_54342;
  wire net_54343;
  wire net_54344;
  wire net_54345;
  wire net_54348;
  wire net_54349;
  wire net_54356;
  wire net_54363;
  wire net_54369;
  wire net_54372;
  wire net_54373;
  wire net_54374;
  wire net_54375;
  wire net_54376;
  wire net_54377;
  wire net_54379;
  wire net_54380;
  wire net_54381;
  wire net_54382;
  wire net_54383;
  wire net_54384;
  wire net_54385;
  wire net_54386;
  wire net_54395;
  wire net_54397;
  wire net_54406;
  wire net_54407;
  wire net_54409;
  wire net_54412;
  wire net_54414;
  wire net_54426;
  wire net_54427;
  wire net_54428;
  wire net_54431;
  wire net_54433;
  wire net_54434;
  wire net_54435;
  wire net_54437;
  wire net_54442;
  wire net_54444;
  wire net_54446;
  wire net_54447;
  wire net_54449;
  wire net_54450;
  wire net_54451;
  wire net_54453;
  wire net_54454;
  wire net_54455;
  wire net_54456;
  wire net_54459;
  wire net_54461;
  wire net_54467;
  wire net_54471;
  wire net_54472;
  wire net_54473;
  wire net_54474;
  wire net_54478;
  wire net_54480;
  wire net_54483;
  wire net_54489;
  wire net_54490;
  wire net_54491;
  wire net_54492;
  wire net_54496;
  wire net_54499;
  wire net_54500;
  wire net_54502;
  wire net_54503;
  wire net_54504;
  wire net_54505;
  wire net_54506;
  wire net_54507;
  wire net_54508;
  wire net_54509;
  wire net_54514;
  wire net_54519;
  wire net_54525;
  wire net_54527;
  wire net_54536;
  wire net_54537;
  wire net_54545;
  wire net_54548;
  wire net_54553;
  wire net_54555;
  wire net_54559;
  wire net_54560;
  wire net_54561;
  wire net_54562;
  wire net_54564;
  wire net_54565;
  wire net_54569;
  wire net_54570;
  wire net_54572;
  wire net_54573;
  wire net_54576;
  wire net_54577;
  wire net_54578;
  wire net_54579;
  wire net_54582;
  wire net_54589;
  wire net_54595;
  wire net_54596;
  wire net_54603;
  wire net_54609;
  wire net_54614;
  wire net_54618;
  wire net_54619;
  wire net_54620;
  wire net_54621;
  wire net_54622;
  wire net_54623;
  wire net_54625;
  wire net_54626;
  wire net_54628;
  wire net_54629;
  wire net_54630;
  wire net_54631;
  wire net_54632;
  wire net_54637;
  wire net_54641;
  wire net_54642;
  wire net_54652;
  wire net_54668;
  wire net_54670;
  wire net_54672;
  wire net_54677;
  wire net_54680;
  wire net_54682;
  wire net_54685;
  wire net_54686;
  wire net_54687;
  wire net_54689;
  wire net_54690;
  wire net_54692;
  wire net_54693;
  wire net_54694;
  wire net_54695;
  wire net_54696;
  wire net_54697;
  wire net_54698;
  wire net_54700;
  wire net_54701;
  wire net_54704;
  wire net_54706;
  wire net_54707;
  wire net_54708;
  wire net_54710;
  wire net_54712;
  wire net_54713;
  wire net_54714;
  wire net_54716;
  wire net_54718;
  wire net_54719;
  wire net_54720;
  wire net_54722;
  wire net_54724;
  wire net_54725;
  wire net_54726;
  wire net_54728;
  wire net_54730;
  wire net_54731;
  wire net_54732;
  wire net_54734;
  wire net_54736;
  wire net_54737;
  wire net_54738;
  wire net_54740;
  wire net_54742;
  wire net_54743;
  wire net_54744;
  wire net_54745;
  wire net_54746;
  wire net_54749;
  wire net_54750;
  wire net_54751;
  wire net_54753;
  wire net_54755;
  wire net_54764;
  wire net_54777;
  wire net_54784;
  wire net_54789;
  wire net_54792;
  wire net_54793;
  wire net_54795;
  wire net_54797;
  wire net_54801;
  wire net_54803;
  wire net_54805;
  wire net_54806;
  wire net_54808;
  wire net_54811;
  wire net_54812;
  wire net_54814;
  wire net_54815;
  wire net_54816;
  wire net_54818;
  wire net_54820;
  wire net_54821;
  wire net_54823;
  wire net_54824;
  wire net_54825;
  wire net_54827;
  wire net_54829;
  wire net_54830;
  wire net_54831;
  wire net_54833;
  wire net_54835;
  wire net_54836;
  wire net_54837;
  wire net_54839;
  wire net_54841;
  wire net_54842;
  wire net_54843;
  wire net_54845;
  wire net_54847;
  wire net_54848;
  wire net_54849;
  wire net_54851;
  wire net_54853;
  wire net_54854;
  wire net_54855;
  wire net_54857;
  wire net_54859;
  wire net_54860;
  wire net_54861;
  wire net_54865;
  wire net_54866;
  wire net_54867;
  wire net_54868;
  wire net_54869;
  wire net_54871;
  wire net_54872;
  wire net_54874;
  wire net_54875;
  wire net_54876;
  wire net_54878;
  wire net_54889;
  wire net_54900;
  wire net_54912;
  wire net_54933;
  wire net_54943;
  wire net_54964;
  wire net_54970;
  wire net_54976;
  wire net_54991;
  wire net_54992;
  wire net_54994;
  wire net_54995;
  wire net_55000;
  wire net_55001;
  wire net_55011;
  wire net_55018;
  wire net_55020;
  wire net_55042;
  wire net_55043;
  wire net_55049;
  wire net_55050;
  wire net_55052;
  wire net_55053;
  wire net_55055;
  wire net_55056;
  wire net_55057;
  wire net_55058;
  wire net_55062;
  wire net_55063;
  wire net_55064;
  wire net_55066;
  wire net_55074;
  wire net_55075;
  wire net_55076;
  wire net_55077;
  wire net_55082;
  wire net_55092;
  wire net_55093;
  wire net_55094;
  wire net_55095;
  wire net_55104;
  wire net_55105;
  wire net_55106;
  wire net_55107;
  wire net_55112;
  wire net_55114;
  wire net_55115;
  wire net_55117;
  wire net_55118;
  wire net_55119;
  wire net_55121;
  wire net_55122;
  wire net_55124;
  wire net_55128;
  wire net_55133;
  wire net_55139;
  wire net_55169;
  wire net_55171;
  wire net_55172;
  wire net_55175;
  wire net_55176;
  wire net_55178;
  wire net_55181;
  wire net_55182;
  wire net_55183;
  wire net_55186;
  wire net_55187;
  wire net_55189;
  wire net_55194;
  wire net_55200;
  wire net_55212;
  wire net_55217;
  wire net_55223;
  wire net_55227;
  wire net_55228;
  wire net_55229;
  wire net_55230;
  wire net_55233;
  wire net_55234;
  wire net_55235;
  wire net_55236;
  wire net_55237;
  wire net_55238;
  wire net_55247;
  wire net_55250;
  wire net_55260;
  wire net_55309;
  wire net_55351;
  wire net_55381;
  wire net_55405;
  wire net_55417;
  wire net_55418;
  wire net_55422;
  wire net_55423;
  wire net_55433;
  wire net_55443;
  wire net_55455;
  wire net_55456;
  wire net_55457;
  wire net_55458;
  wire net_55470;
  wire net_55479;
  wire net_55480;
  wire net_55481;
  wire net_55482;
  wire net_55483;
  wire net_55484;
  wire net_55858;
  wire net_55859;
  wire net_55880;
  wire net_55979;
  wire net_55980;
  wire net_55983;
  wire net_56021;
  wire net_56024;
  wire net_56025;
  wire net_56026;
  wire net_56030;
  wire net_56031;
  wire net_56034;
  wire net_56036;
  wire net_56037;
  wire net_56040;
  wire net_56047;
  wire net_56064;
  wire net_56065;
  wire net_56066;
  wire net_56067;
  wire net_56076;
  wire net_56079;
  wire net_56082;
  wire net_56084;
  wire net_56085;
  wire net_56088;
  wire net_56089;
  wire net_56090;
  wire net_56091;
  wire net_56094;
  wire net_56095;
  wire net_56098;
  wire net_56099;
  wire net_56102;
  wire net_56244;
  wire net_56245;
  wire net_56515;
  wire net_56521;
  wire net_56522;
  wire net_56523;
  wire net_56534;
  wire net_56535;
  wire net_56584;
  wire net_56697;
  wire net_56698;
  wire net_56699;
  wire net_56700;
  wire net_56703;
  wire net_56732;
  wire net_56776;
  wire net_56777;
  wire net_56780;
  wire net_56785;
  wire net_56790;
  wire net_56793;
  wire net_56800;
  wire net_56805;
  wire net_56819;
  wire net_56821;
  wire net_56825;
  wire net_56826;
  wire net_56827;
  wire net_56828;
  wire net_56838;
  wire net_56839;
  wire net_56840;
  wire net_56843;
  wire net_56844;
  wire net_56845;
  wire net_56846;
  wire net_56857;
  wire net_56858;
  wire net_56859;
  wire net_56860;
  wire net_56861;
  wire net_56862;
  wire net_56863;
  wire net_56870;
  wire net_56897;
  wire net_56898;
  wire net_56899;
  wire net_56904;
  wire net_56905;
  wire net_56906;
  wire net_56908;
  wire net_56909;
  wire net_56911;
  wire net_56912;
  wire net_56914;
  wire net_56915;
  wire net_56916;
  wire net_56917;
  wire net_56920;
  wire net_56921;
  wire net_56924;
  wire net_56928;
  wire net_56930;
  wire net_56931;
  wire net_56932;
  wire net_56933;
  wire net_56937;
  wire net_56938;
  wire net_56939;
  wire net_56942;
  wire net_56943;
  wire net_56948;
  wire net_56949;
  wire net_56950;
  wire net_56951;
  wire net_56954;
  wire net_56955;
  wire net_56956;
  wire net_56957;
  wire net_56960;
  wire net_56961;
  wire net_56962;
  wire net_56963;
  wire net_56966;
  wire net_56967;
  wire net_56968;
  wire net_56969;
  wire net_56972;
  wire net_56976;
  wire net_56977;
  wire net_57023;
  wire net_57027;
  wire net_57028;
  wire net_57030;
  wire net_57034;
  wire net_57038;
  wire net_57041;
  wire net_57044;
  wire net_57046;
  wire net_57049;
  wire net_57051;
  wire net_57053;
  wire net_57054;
  wire net_57056;
  wire net_57059;
  wire net_57061;
  wire net_57066;
  wire net_57068;
  wire net_57078;
  wire net_57080;
  wire net_57083;
  wire net_57085;
  wire net_57097;
  wire net_57098;
  wire net_57099;
  wire net_57100;
  wire net_57227;
  wire net_57259;
  wire net_57391;
  wire net_57403;
  wire net_57410;
  wire net_57412;
  wire net_57414;
  wire net_57415;
  wire net_57418;
  wire net_57428;
  wire net_57430;
  wire net_57458;
  wire net_57459;
  wire net_57460;
  wire net_57461;
  wire net_57464;
  wire net_57466;
  wire net_57468;
  wire net_57469;
  wire net_57471;
  wire net_57495;
  wire net_57515;
  wire net_57518;
  wire net_57523;
  wire net_57526;
  wire net_57527;
  wire net_57528;
  wire net_57529;
  wire net_57535;
  wire net_57536;
  wire net_57539;
  wire net_57541;
  wire net_57543;
  wire net_57569;
  wire net_57570;
  wire net_57571;
  wire net_57572;
  wire net_57575;
  wire net_57576;
  wire net_57578;
  wire net_57581;
  wire net_57582;
  wire net_57583;
  wire net_57584;
  wire net_57587;
  wire net_57588;
  wire net_57589;
  wire net_57590;
  wire net_57591;
  wire net_57592;
  wire net_57594;
  wire net_57599;
  wire net_57601;
  wire net_57616;
  wire net_57625;
  wire net_57635;
  wire net_57636;
  wire net_57640;
  wire net_57641;
  wire net_57642;
  wire net_57643;
  wire net_57647;
  wire net_57649;
  wire net_57652;
  wire net_57660;
  wire net_57669;
  wire net_57673;
  wire net_57675;
  wire net_57676;
  wire net_57679;
  wire net_57681;
  wire net_57682;
  wire net_57683;
  wire net_57685;
  wire net_57687;
  wire net_57688;
  wire net_57689;
  wire net_57691;
  wire net_57693;
  wire net_57694;
  wire net_57695;
  wire net_57697;
  wire net_57699;
  wire net_57700;
  wire net_57701;
  wire net_57703;
  wire net_57705;
  wire net_57706;
  wire net_57707;
  wire net_57710;
  wire net_57712;
  wire net_57713;
  wire net_57719;
  wire net_57721;
  wire net_57722;
  wire net_57723;
  wire net_57742;
  wire net_57751;
  wire net_57763;
  wire net_57764;
  wire net_57776;
  wire net_57779;
  wire net_57833;
  wire net_57834;
  wire net_57835;
  wire net_57836;
  wire net_57841;
  wire net_57842;
  wire net_57843;
  wire net_57844;
  wire net_57845;
  wire net_57846;
  wire net_57847;
  wire net_57863;
  wire net_57867;
  wire net_57868;
  wire net_57870;
  wire net_57884;
  wire net_57885;
  wire net_57887;
  wire net_57888;
  wire net_57890;
  wire net_57893;
  wire net_57897;
  wire net_57899;
  wire net_57900;
  wire net_57902;
  wire net_57903;
  wire net_57915;
  wire net_57920;
  wire net_57926;
  wire net_57927;
  wire net_57928;
  wire net_57929;
  wire net_57933;
  wire net_57938;
  wire net_57939;
  wire net_57940;
  wire net_57941;
  wire net_57944;
  wire net_57952;
  wire net_57959;
  wire net_57960;
  wire net_57961;
  wire net_57963;
  wire net_57964;
  wire net_57965;
  wire net_57966;
  wire net_57967;
  wire net_57968;
  wire net_57969;
  wire net_57970;
  wire net_57978;
  wire net_57981;
  wire net_57988;
  wire net_57992;
  wire net_57993;
  wire net_57995;
  wire net_58006;
  wire net_58007;
  wire net_58012;
  wire net_58013;
  wire net_58014;
  wire net_58015;
  wire net_58018;
  wire net_58019;
  wire net_58021;
  wire net_58023;
  wire net_58024;
  wire net_58026;
  wire net_58027;
  wire net_58031;
  wire net_58034;
  wire net_58035;
  wire net_58037;
  wire net_58038;
  wire net_58039;
  wire net_58040;
  wire net_58043;
  wire net_58049;
  wire net_58050;
  wire net_58051;
  wire net_58052;
  wire net_58055;
  wire net_58056;
  wire net_58057;
  wire net_58058;
  wire net_58064;
  wire net_58067;
  wire net_58076;
  wire net_58079;
  wire net_58080;
  wire net_58081;
  wire net_58082;
  wire net_58083;
  wire net_58084;
  wire net_58086;
  wire net_58087;
  wire net_58088;
  wire net_58089;
  wire net_58090;
  wire net_58091;
  wire net_58092;
  wire net_58093;
  wire net_58102;
  wire net_58110;
  wire net_58121;
  wire net_58128;
  wire net_58129;
  wire net_58130;
  wire net_58133;
  wire net_58134;
  wire net_58135;
  wire net_58136;
  wire net_58137;
  wire net_58138;
  wire net_58140;
  wire net_58141;
  wire net_58142;
  wire net_58144;
  wire net_58145;
  wire net_58147;
  wire net_58148;
  wire net_58149;
  wire net_58150;
  wire net_58151;
  wire net_58152;
  wire net_58154;
  wire net_58155;
  wire net_58156;
  wire net_58157;
  wire net_58158;
  wire net_58160;
  wire net_58166;
  wire net_58167;
  wire net_58168;
  wire net_58169;
  wire net_58172;
  wire net_58173;
  wire net_58174;
  wire net_58175;
  wire net_58178;
  wire net_58179;
  wire net_58180;
  wire net_58181;
  wire net_58184;
  wire net_58185;
  wire net_58186;
  wire net_58187;
  wire net_58190;
  wire net_58191;
  wire net_58192;
  wire net_58193;
  wire net_58196;
  wire net_58197;
  wire net_58198;
  wire net_58199;
  wire net_58203;
  wire net_58206;
  wire net_58207;
  wire net_58209;
  wire net_58210;
  wire net_58211;
  wire net_58212;
  wire net_58213;
  wire net_58214;
  wire net_58215;
  wire net_58216;
  wire net_58222;
  wire net_58223;
  wire net_58225;
  wire net_58229;
  wire net_58230;
  wire net_58231;
  wire net_58234;
  wire net_58236;
  wire net_58240;
  wire net_58241;
  wire net_58243;
  wire net_58244;
  wire net_58258;
  wire net_58260;
  wire net_58261;
  wire net_58262;
  wire net_58263;
  wire net_58264;
  wire net_58270;
  wire net_58272;
  wire net_58273;
  wire net_58274;
  wire net_58276;
  wire net_58277;
  wire net_58279;
  wire net_58280;
  wire net_58281;
  wire net_58283;
  wire net_58284;
  wire net_58285;
  wire net_58286;
  wire net_58290;
  wire net_58291;
  wire net_58295;
  wire net_58296;
  wire net_58297;
  wire net_58298;
  wire net_58302;
  wire net_58309;
  wire net_58310;
  wire net_58315;
  wire net_58319;
  wire net_58325;
  wire net_58326;
  wire net_58327;
  wire net_58328;
  wire net_58329;
  wire net_58330;
  wire net_58332;
  wire net_58333;
  wire net_58334;
  wire net_58335;
  wire net_58336;
  wire net_58337;
  wire net_58338;
  wire net_58339;
  wire net_58344;
  wire net_58349;
  wire net_58358;
  wire net_58359;
  wire net_58367;
  wire net_58382;
  wire net_58383;
  wire net_58386;
  wire net_58387;
  wire net_58391;
  wire net_58392;
  wire net_58395;
  wire net_58396;
  wire net_58397;
  wire net_58398;
  wire net_58402;
  wire net_58403;
  wire net_58404;
  wire net_58407;
  wire net_58414;
  wire net_58415;
  wire net_58420;
  wire net_58424;
  wire net_58425;
  wire net_58426;
  wire net_58427;
  wire net_58432;
  wire net_58437;
  wire net_58438;
  wire net_58445;
  wire net_58448;
  wire net_58452;
  wire net_58453;
  wire net_58455;
  wire net_58458;
  wire net_58459;
  wire net_58460;
  wire net_58461;
  wire net_58462;
  wire net_58489;
  wire net_58498;
  wire net_58500;
  wire net_58501;
  wire net_58504;
  wire net_58509;
  wire net_58511;
  wire net_58513;
  wire net_58517;
  wire net_58518;
  wire net_58520;
  wire net_58521;
  wire net_58523;
  wire net_58531;
  wire net_58535;
  wire net_58536;
  wire net_58537;
  wire net_58538;
  wire net_58550;
  wire net_58553;
  wire net_58555;
  wire net_58559;
  wire net_58568;
  wire net_58571;
  wire net_58575;
  wire net_58576;
  wire net_58578;
  wire net_58579;
  wire net_58580;
  wire net_58581;
  wire net_58583;
  wire net_58584;
  wire net_58585;
  wire net_58609;
  wire net_58620;
  wire net_58630;
  wire net_58633;
  wire net_58644;
  wire net_58645;
  wire net_58650;
  wire net_58658;
  wire net_58665;
  wire net_58671;
  wire net_58682;
  wire net_58685;
  wire net_58695;
  wire net_58698;
  wire net_58699;
  wire net_58701;
  wire net_58702;
  wire net_58703;
  wire net_58705;
  wire net_58707;
  wire net_58708;
  wire net_58726;
  wire net_58735;
  wire net_58745;
  wire net_58747;
  wire net_58749;
  wire net_58753;
  wire net_58758;
  wire net_58759;
  wire net_58760;
  wire net_58761;
  wire net_58763;
  wire net_58764;
  wire net_58766;
  wire net_58767;
  wire net_58769;
  wire net_58776;
  wire net_58778;
  wire net_58781;
  wire net_58793;
  wire net_58796;
  wire net_58799;
  wire net_58800;
  wire net_58801;
  wire net_58802;
  wire net_58808;
  wire net_58817;
  wire net_58818;
  wire net_58819;
  wire net_58820;
  wire net_58821;
  wire net_58822;
  wire net_58824;
  wire net_58827;
  wire net_58829;
  wire net_58830;
  wire net_58837;
  wire net_58846;
  wire net_58847;
  wire net_58850;
  wire net_58852;
  wire net_58853;
  wire net_58865;
  wire net_58867;
  wire net_58873;
  wire net_58875;
  wire net_58877;
  wire net_58884;
  wire net_58892;
  wire net_58894;
  wire net_58899;
  wire net_58904;
  wire net_58905;
  wire net_58906;
  wire net_58907;
  wire net_58935;
  wire net_58936;
  wire net_58941;
  wire net_58943;
  wire net_58944;
  wire net_58945;
  wire net_58947;
  wire net_58949;
  wire net_58953;
  wire net_58954;
  wire net_58962;
  wire net_58971;
  wire net_58973;
  wire net_58980;
  wire net_58988;
  wire net_58990;
  wire net_58991;
  wire net_58992;
  wire net_58993;
  wire net_58994;
  wire net_58995;
  wire net_58999;
  wire net_59002;
  wire net_59004;
  wire net_59005;
  wire net_59014;
  wire net_59016;
  wire net_59017;
  wire net_59023;
  wire net_59027;
  wire net_59029;
  wire net_59035;
  wire net_59046;
  wire net_59051;
  wire net_59052;
  wire net_59053;
  wire net_59054;
  wire net_59063;
  wire net_59064;
  wire net_59065;
  wire net_59066;
  wire net_59067;
  wire net_59068;
  wire net_59076;
  wire net_59084;
  wire net_59105;
  wire net_59140;
  wire net_59187;
  wire net_59190;
  wire net_59191;
  wire net_59197;
  wire net_59198;
  wire net_59206;
  wire net_59218;
  wire net_59219;
  wire net_59317;
  wire net_59321;
  wire net_59323;
  wire net_59351;
  wire net_59567;
  wire net_59589;
  wire net_59597;
  wire net_59709;
  wire net_59735;
  wire net_59737;
  wire net_59753;
  wire net_59778;
  wire net_59783;
  wire net_59785;
  wire net_59805;
  wire net_59806;
  wire net_59813;
  wire net_59838;
  wire net_59842;
  wire net_59851;
  wire net_59859;
  wire net_59862;
  wire net_59867;
  wire net_59869;
  wire net_59870;
  wire net_59875;
  wire net_59879;
  wire net_59888;
  wire net_59889;
  wire net_59890;
  wire net_59891;
  wire net_59895;
  wire net_59913;
  wire net_59914;
  wire net_59915;
  wire net_59928;
  wire net_59929;
  wire net_59931;
  wire net_59932;
  wire net_59935;
  wire net_59936;
  wire net_59938;
  wire net_59984;
  wire net_59988;
  wire net_60011;
  wire net_60014;
  wire net_60059;
  wire net_60061;
  wire net_60528;
  wire net_60529;
  wire net_60530;
  wire net_60532;
  wire net_60604;
  wire net_60606;
  wire net_60610;
  wire net_60611;
  wire net_60614;
  wire net_60615;
  wire net_60628;
  wire net_60637;
  wire net_60638;
  wire net_60639;
  wire net_60643;
  wire net_60644;
  wire net_60645;
  wire net_60646;
  wire net_60649;
  wire net_60650;
  wire net_60651;
  wire net_60652;
  wire net_60655;
  wire net_60656;
  wire net_60657;
  wire net_60658;
  wire net_60673;
  wire net_60676;
  wire net_60683;
  wire net_60684;
  wire net_60710;
  wire net_60729;
  wire net_60732;
  wire net_60735;
  wire net_60736;
  wire net_60738;
  wire net_60739;
  wire net_60740;
  wire net_60747;
  wire net_60749;
  wire net_60753;
  wire net_60754;
  wire net_60758;
  wire net_60767;
  wire net_60768;
  wire net_60769;
  wire net_60772;
  wire net_60773;
  wire net_60778;
  wire net_60779;
  wire net_60781;
  wire net_60784;
  wire net_60785;
  wire net_60786;
  wire net_60787;
  wire net_60791;
  wire net_60792;
  wire net_60793;
  wire net_60796;
  wire net_60797;
  wire net_60798;
  wire net_60799;
  wire net_60802;
  wire net_60803;
  wire net_60804;
  wire net_60805;
  wire net_60806;
  wire net_60807;
  wire net_60840;
  wire net_60934;
  wire net_60935;
  wire net_60936;
  wire net_60937;
  wire net_60938;
  wire net_60939;
  wire net_60942;
  wire net_60943;
  wire net_60965;
  wire net_61055;
  wire net_61076;
  wire net_61119;
  wire net_61123;
  wire net_61144;
  wire net_61175;
  wire net_61176;
  wire net_61201;
  wire net_61203;
  wire net_61207;
  wire net_61333;
  wire net_61350;
  wire net_61353;
  wire net_61376;
  wire net_61421;
  wire net_61422;
  wire net_61426;
  wire net_61427;
  wire net_61428;
  wire net_61429;
  wire net_61430;
  wire net_61431;
  wire net_61435;
  wire net_61473;
  wire net_61476;
  wire net_61483;
  wire net_61485;
  wire net_61486;
  wire net_61498;
  wire net_61501;
  wire net_61530;
  wire net_61540;
  wire net_61542;
  wire net_61544;
  wire net_61545;
  wire net_61546;
  wire net_61552;
  wire net_61571;
  wire net_61579;
  wire net_61588;
  wire net_61591;
  wire net_61592;
  wire net_61594;
  wire net_61596;
  wire net_61598;
  wire net_61599;
  wire net_61600;
  wire net_61601;
  wire net_61602;
  wire net_61609;
  wire net_61610;
  wire net_61613;
  wire net_61616;
  wire net_61617;
  wire net_61623;
  wire net_61626;
  wire net_61629;
  wire net_61634;
  wire net_61636;
  wire net_61645;
  wire net_61646;
  wire net_61647;
  wire net_61648;
  wire net_61651;
  wire net_61652;
  wire net_61653;
  wire net_61654;
  wire net_61657;
  wire net_61658;
  wire net_61659;
  wire net_61667;
  wire net_61668;
  wire net_61670;
  wire net_61671;
  wire net_61674;
  wire net_61675;
  wire net_61687;
  wire net_61692;
  wire net_61696;
  wire net_61699;
  wire net_61715;
  wire net_61716;
  wire net_61717;
  wire net_61719;
  wire net_61724;
  wire net_61726;
  wire net_61728;
  wire net_61729;
  wire net_61730;
  wire net_61731;
  wire net_61735;
  wire net_61736;
  wire net_61737;
  wire net_61738;
  wire net_61739;
  wire net_61740;
  wire net_61741;
  wire net_61743;
  wire net_61745;
  wire net_61746;
  wire net_61749;
  wire net_61751;
  wire net_61752;
  wire net_61753;
  wire net_61755;
  wire net_61757;
  wire net_61758;
  wire net_61759;
  wire net_61761;
  wire net_61763;
  wire net_61764;
  wire net_61765;
  wire net_61767;
  wire net_61769;
  wire net_61770;
  wire net_61771;
  wire net_61773;
  wire net_61775;
  wire net_61776;
  wire net_61777;
  wire net_61779;
  wire net_61781;
  wire net_61782;
  wire net_61783;
  wire net_61785;
  wire net_61787;
  wire net_61788;
  wire net_61789;
  wire net_61790;
  wire net_61791;
  wire net_61793;
  wire net_61794;
  wire net_61795;
  wire net_61797;
  wire net_61798;
  wire net_61799;
  wire net_61818;
  wire net_61823;
  wire net_61824;
  wire net_61826;
  wire net_61829;
  wire net_61837;
  wire net_61838;
  wire net_61841;
  wire net_61842;
  wire net_61845;
  wire net_61850;
  wire net_61851;
  wire net_61852;
  wire net_61854;
  wire net_61855;
  wire net_61856;
  wire net_61857;
  wire net_61860;
  wire net_61861;
  wire net_61862;
  wire net_61863;
  wire net_61864;
  wire net_61866;
  wire net_61868;
  wire net_61869;
  wire net_61870;
  wire net_61872;
  wire net_61874;
  wire net_61875;
  wire net_61876;
  wire net_61878;
  wire net_61880;
  wire net_61881;
  wire net_61882;
  wire net_61884;
  wire net_61886;
  wire net_61887;
  wire net_61888;
  wire net_61890;
  wire net_61892;
  wire net_61893;
  wire net_61894;
  wire net_61896;
  wire net_61898;
  wire net_61899;
  wire net_61900;
  wire net_61902;
  wire net_61904;
  wire net_61905;
  wire net_61906;
  wire net_61909;
  wire net_61911;
  wire net_61912;
  wire net_61913;
  wire net_61914;
  wire net_61916;
  wire net_61918;
  wire net_61919;
  wire net_61920;
  wire net_61929;
  wire net_61942;
  wire net_61943;
  wire net_61946;
  wire net_61947;
  wire net_61949;
  wire net_61957;
  wire net_61961;
  wire net_61962;
  wire net_61963;
  wire net_61965;
  wire net_61966;
  wire net_61967;
  wire net_61968;
  wire net_61969;
  wire net_61970;
  wire net_61972;
  wire net_61973;
  wire net_61974;
  wire net_61976;
  wire net_61977;
  wire net_61978;
  wire net_61983;
  wire net_61984;
  wire net_61985;
  wire net_61986;
  wire net_61990;
  wire net_61991;
  wire net_61992;
  wire net_61993;
  wire net_61996;
  wire net_61997;
  wire net_61998;
  wire net_61999;
  wire net_62002;
  wire net_62003;
  wire net_62004;
  wire net_62005;
  wire net_62010;
  wire net_62017;
  wire net_62020;
  wire net_62021;
  wire net_62022;
  wire net_62023;
  wire net_62026;
  wire net_62027;
  wire net_62028;
  wire net_62029;
  wire net_62033;
  wire net_62034;
  wire net_62040;
  wire net_62044;
  wire net_62046;
  wire net_62051;
  wire net_62053;
  wire net_62057;
  wire net_62064;
  wire net_62066;
  wire net_62071;
  wire net_62081;
  wire net_62082;
  wire net_62083;
  wire net_62086;
  wire net_62089;
  wire net_62090;
  wire net_62092;
  wire net_62094;
  wire net_62095;
  wire net_62096;
  wire net_62098;
  wire net_62100;
  wire net_62101;
  wire net_62105;
  wire net_62111;
  wire net_62116;
  wire net_62119;
  wire net_62120;
  wire net_62121;
  wire net_62122;
  wire net_62125;
  wire net_62132;
  wire net_62137;
  wire net_62138;
  wire net_62139;
  wire net_62140;
  wire net_62145;
  wire net_62149;
  wire net_62155;
  wire net_62156;
  wire net_62157;
  wire net_62158;
  wire net_62159;
  wire net_62160;
  wire net_62162;
  wire net_62164;
  wire net_62165;
  wire net_62166;
  wire net_62167;
  wire net_62168;
  wire net_62169;
  wire net_62178;
  wire net_62184;
  wire net_62189;
  wire net_62204;
  wire net_62206;
  wire net_62208;
  wire net_62209;
  wire net_62210;
  wire net_62217;
  wire net_62218;
  wire net_62220;
  wire net_62221;
  wire net_62224;
  wire net_62227;
  wire net_62229;
  wire net_62230;
  wire net_62232;
  wire net_62239;
  wire net_62243;
  wire net_62248;
  wire net_62249;
  wire net_62250;
  wire net_62251;
  wire net_62256;
  wire net_62260;
  wire net_62261;
  wire net_62262;
  wire net_62263;
  wire net_62266;
  wire net_62268;
  wire net_62275;
  wire net_62280;
  wire net_62282;
  wire net_62283;
  wire net_62286;
  wire net_62287;
  wire net_62298;
  wire net_62303;
  wire net_62304;
  wire net_62307;
  wire net_62308;
  wire net_62320;
  wire net_62327;
  wire net_62331;
  wire net_62334;
  wire net_62337;
  wire net_62339;
  wire net_62340;
  wire net_62344;
  wire net_62346;
  wire net_62348;
  wire net_62350;
  wire net_62353;
  wire net_62354;
  wire net_62356;
  wire net_62359;
  wire net_62360;
  wire net_62377;
  wire net_62378;
  wire net_62383;
  wire net_62384;
  wire net_62385;
  wire net_62386;
  wire net_62392;
  wire net_62395;
  wire net_62396;
  wire net_62398;
  wire net_62402;
  wire net_62403;
  wire net_62405;
  wire net_62406;
  wire net_62409;
  wire net_62428;
  wire net_62438;
  wire net_62456;
  wire net_62457;
  wire net_62458;
  wire net_62460;
  wire net_62467;
  wire net_62469;
  wire net_62470;
  wire net_62471;
  wire net_62472;
  wire net_62478;
  wire net_62479;
  wire net_62484;
  wire net_62488;
  wire net_62489;
  wire net_62490;
  wire net_62491;
  wire net_62495;
  wire net_62502;
  wire net_62503;
  wire net_62513;
  wire net_62515;
  wire net_62519;
  wire net_62526;
  wire net_62528;
  wire net_62529;
  wire net_62533;
  wire net_62534;
  wire net_62535;
  wire net_62548;
  wire net_62555;
  wire net_62566;
  wire net_62572;
  wire net_62573;
  wire net_62574;
  wire net_62578;
  wire net_62579;
  wire net_62582;
  wire net_62584;
  wire net_62588;
  wire net_62589;
  wire net_62592;
  wire net_62593;
  wire net_62597;
  wire net_62599;
  wire net_62600;
  wire net_62605;
  wire net_62606;
  wire net_62607;
  wire net_62608;
  wire net_62611;
  wire net_62612;
  wire net_62613;
  wire net_62614;
  wire net_62619;
  wire net_62632;
  wire net_62641;
  wire net_62642;
  wire net_62643;
  wire net_62644;
  wire net_62650;
  wire net_62651;
  wire net_62652;
  wire net_62655;
  wire net_62657;
  wire net_62658;
  wire net_62659;
  wire net_62660;
  wire net_62661;
  wire net_62662;
  wire net_62666;
  wire net_62702;
  wire net_62703;
  wire net_62706;
  wire net_62715;
  wire net_62720;
  wire net_62722;
  wire net_62723;
  wire net_62724;
  wire net_62729;
  wire net_62746;
  wire net_62747;
  wire net_62748;
  wire net_62761;
  wire net_62764;
  wire net_62766;
  wire net_62774;
  wire net_62775;
  wire net_62778;
  wire net_62779;
  wire net_62780;
  wire net_62781;
  wire net_62782;
  wire net_62784;
  wire net_62789;
  wire net_62797;
  wire net_62802;
  wire net_62818;
  wire net_62821;
  wire net_62828;
  wire net_62829;
  wire net_62833;
  wire net_62834;
  wire net_62838;
  wire net_62844;
  wire net_62849;
  wire net_62851;
  wire net_62863;
  wire net_62865;
  wire net_62887;
  wire net_62888;
  wire net_62889;
  wire net_62890;
  wire net_62894;
  wire net_62895;
  wire net_62897;
  wire net_62898;
  wire net_62899;
  wire net_62907;
  wire net_62956;
  wire net_62967;
  wire net_63010;
  wire net_63011;
  wire net_63068;
  wire net_63079;
  wire net_63091;
  wire net_63121;
  wire net_63130;
  wire net_63143;
  wire net_63144;
  wire net_63180;
  wire net_63191;
  wire net_63192;
  wire net_63200;
  wire net_63204;
  wire net_63205;
  wire net_63228;
  wire net_63250;
  wire net_63251;
  wire net_63252;
  wire net_63253;
  wire net_63262;
  wire net_63263;
  wire net_63264;
  wire net_63265;
  wire net_63266;
  wire net_63267;
  wire net_63418;
  wire net_63439;
  wire net_63444;
  wire net_63499;
  wire net_63512;
  wire net_63513;
  wire net_63548;
  wire net_63683;
  wire net_63710;
  wire net_63743;
  wire net_63745;
  wire net_63762;
  wire net_63763;
  wire net_63764;
  wire net_63765;
  wire net_63766;
  wire net_63767;
  wire net_63768;
  wire net_63807;
  wire net_63819;
  wire net_63823;
  wire net_63824;
  wire net_63829;
  wire net_63830;
  wire net_63831;
  wire net_63835;
  wire net_63836;
  wire net_63837;
  wire net_63838;
  wire net_63841;
  wire net_63842;
  wire net_63859;
  wire net_63860;
  wire net_63861;
  wire net_63862;
  wire net_63865;
  wire net_63866;
  wire net_63867;
  wire net_63868;
  wire net_63877;
  wire net_63878;
  wire net_63879;
  wire net_63880;
  wire net_63884;
  wire net_63886;
  wire net_63888;
  wire net_63890;
  wire net_63914;
  wire net_63928;
  wire net_63930;
  wire net_63934;
  wire net_63936;
  wire net_63938;
  wire net_63939;
  wire net_63954;
  wire net_63988;
  wire net_63989;
  wire net_63990;
  wire net_63991;
  wire net_64001;
  wire net_64002;
  wire net_64003;
  wire net_64354;
  wire net_64355;
  wire net_64390;
  wire net_64392;
  wire net_64410;
  wire net_64436;
  wire net_64443;
  wire net_64444;
  wire net_64449;
  wire net_64455;
  wire net_64458;
  wire net_64461;
  wire net_64462;
  wire net_64466;
  wire net_64475;
  wire net_64480;
  wire net_64481;
  wire net_64483;
  wire net_64486;
  wire net_64488;
  wire net_64498;
  wire net_64499;
  wire net_64500;
  wire net_64501;
  wire net_64514;
  wire net_64515;
  wire net_64763;
  wire net_64764;
  wire net_64765;
  wire net_64766;
  wire net_64768;
  wire net_64769;
  wire net_64770;
  wire net_64773;
  wire net_64814;
  wire net_64818;
  wire net_64820;
  wire net_64827;
  wire net_64829;
  wire net_64830;
  wire net_64831;
  wire net_64834;
  wire net_64838;
  wire net_64842;
  wire net_64845;
  wire net_64848;
  wire net_64850;
  wire net_64852;
  wire net_64854;
  wire net_64856;
  wire net_64858;
  wire net_64860;
  wire net_64862;
  wire net_64864;
  wire net_64866;
  wire net_64868;
  wire net_64870;
  wire net_64872;
  wire net_64874;
  wire net_64876;
  wire net_64878;
  wire net_64880;
  wire net_64882;
  wire net_64886;
  wire net_64890;
  wire net_64891;
  wire net_64893;
  wire net_64922;
  wire net_64943;
  wire net_64962;
  wire net_64963;
  wire net_65029;
  wire net_65256;
  wire net_65290;
  wire net_65298;
  wire net_65302;
  wire net_65304;
  wire net_65307;
  wire net_65308;
  wire net_65315;
  wire net_65318;
  wire net_65321;
  wire net_65341;
  wire net_65342;
  wire net_65343;
  wire net_65344;
  wire net_65350;
  wire net_65355;
  wire net_65359;
  wire net_65360;
  wire net_65361;
  wire net_65362;
  wire net_65367;
  wire net_65371;
  wire net_65372;
  wire net_65375;
  wire net_65376;
  wire net_65428;
  wire net_65485;
  wire net_65547;
  wire net_65548;
  wire net_65552;
  wire net_65566;
  wire net_65576;
  wire net_65583;
  wire net_65600;
  wire net_65608;
  wire net_65621;
  wire net_65622;
  wire net_65625;
  wire net_65658;
  wire net_65667;
  wire net_65674;
  wire net_65675;
  wire net_65677;
  wire net_65678;
  wire net_65679;
  wire net_65680;
  wire net_65683;
  wire net_65684;
  wire net_65686;
  wire net_65687;
  wire net_65688;
  wire net_65689;
  wire net_65693;
  wire net_65695;
  wire net_65698;
  wire net_65699;
  wire net_65700;
  wire net_65701;
  wire net_65704;
  wire net_65705;
  wire net_65706;
  wire net_65707;
  wire net_65712;
  wire net_65723;
  wire net_65728;
  wire net_65729;
  wire net_65730;
  wire net_65731;
  wire net_65734;
  wire net_65735;
  wire net_65736;
  wire net_65737;
  wire net_65744;
  wire net_65745;
  wire net_65750;
  wire net_65753;
  wire net_65759;
  wire net_65763;
  wire net_65767;
  wire net_65768;
  wire net_65790;
  wire net_65791;
  wire net_65792;
  wire net_65801;
  wire net_65806;
  wire net_65807;
  wire net_65812;
  wire net_65814;
  wire net_65821;
  wire net_65833;
  wire net_65834;
  wire net_65835;
  wire net_65836;
  wire net_65842;
  wire net_65846;
  wire net_65848;
  wire net_65868;
  wire net_65870;
  wire net_65872;
  wire net_65873;
  wire net_65874;
  wire net_65875;
  wire net_65877;
  wire net_65878;
  wire net_65886;
  wire net_65888;
  wire net_65893;
  wire net_65897;
  wire net_65903;
  wire net_65917;
  wire net_65918;
  wire net_65935;
  wire net_65937;
  wire net_65942;
  wire net_65952;
  wire net_65953;
  wire net_65974;
  wire net_65976;
  wire net_65987;
  wire net_65990;
  wire net_65991;
  wire net_65993;
  wire net_65996;
  wire net_65997;
  wire net_66024;
  wire net_66034;
  wire net_66035;
  wire net_66036;
  wire net_66040;
  wire net_66041;
  wire net_66042;
  wire net_66049;
  wire net_66050;
  wire net_66054;
  wire net_66055;
  wire net_66056;
  wire net_66057;
  wire net_66061;
  wire net_66062;
  wire net_66065;
  wire net_66068;
  wire net_66069;
  wire net_66079;
  wire net_66080;
  wire net_66081;
  wire net_66082;
  wire net_66085;
  wire net_66087;
  wire net_66091;
  wire net_66094;
  wire net_66097;
  wire net_66098;
  wire net_66099;
  wire net_66100;
  wire net_66103;
  wire net_66104;
  wire net_66105;
  wire net_66106;
  wire net_66110;
  wire net_66113;
  wire net_66114;
  wire net_66117;
  wire net_66123;
  wire net_66130;
  wire net_66134;
  wire net_66135;
  wire net_66158;
  wire net_66178;
  wire net_66181;
  wire net_66184;
  wire net_66196;
  wire net_66198;
  wire net_66203;
  wire net_66236;
  wire net_66237;
  wire net_66239;
  wire net_66240;
  wire net_66241;
  wire net_66244;
  wire net_66246;
  wire net_66255;
  wire net_66256;
  wire net_66281;
  wire net_66321;
  wire net_66359;
  wire net_66360;
  wire net_66362;
  wire net_66363;
  wire net_66364;
  wire net_66365;
  wire net_66366;
  wire net_66368;
  wire net_66369;
  wire net_66379;
  wire net_66382;
  wire net_66405;
  wire net_66408;
  wire net_66414;
  wire net_66415;
  wire net_66416;
  wire net_66422;
  wire net_66430;
  wire net_66433;
  wire net_66448;
  wire net_66449;
  wire net_66450;
  wire net_66451;
  wire net_66456;
  wire net_66460;
  wire net_66463;
  wire net_66482;
  wire net_66483;
  wire net_66486;
  wire net_66489;
  wire net_66490;
  wire net_66491;
  wire net_66492;
  wire net_66498;
  wire net_66500;
  wire net_66502;
  wire net_66503;
  wire net_66505;
  wire net_66515;
  wire net_66517;
  wire net_66527;
  wire net_66528;
  wire net_66531;
  wire net_66533;
  wire net_66537;
  wire net_66538;
  wire net_66543;
  wire net_66546;
  wire net_66553;
  wire net_66554;
  wire net_66557;
  wire net_66565;
  wire net_66566;
  wire net_66567;
  wire net_66568;
  wire net_66577;
  wire net_66585;
  wire net_66589;
  wire net_66590;
  wire net_66591;
  wire net_66592;
  wire net_66596;
  wire net_66597;
  wire net_66601;
  wire net_66605;
  wire net_66606;
  wire net_66608;
  wire net_66609;
  wire net_66610;
  wire net_66613;
  wire net_66614;
  wire net_66650;
  wire net_66652;
  wire net_66653;
  wire net_66656;
  wire net_66658;
  wire net_66660;
  wire net_66661;
  wire net_66664;
  wire net_66667;
  wire net_66674;
  wire net_66675;
  wire net_66676;
  wire net_66690;
  wire net_66696;
  wire net_66700;
  wire net_66701;
  wire net_66702;
  wire net_66703;
  wire net_66708;
  wire net_66712;
  wire net_66713;
  wire net_66714;
  wire net_66715;
  wire net_66724;
  wire net_66728;
  wire net_66729;
  wire net_66736;
  wire net_66737;
  wire net_66797;
  wire net_66850;
  wire net_66851;
  wire net_66852;
  wire net_67633;
  wire net_67635;
  wire net_67637;
  wire net_67642;
  wire net_67643;
  wire net_67645;
  wire net_67647;
  wire net_67649;
  wire net_67650;
  wire net_67654;
  wire net_67656;
  wire net_67657;
  wire net_67660;
  wire net_67672;
  wire net_67673;
  wire net_67674;
  wire net_67675;
  wire net_67678;
  wire net_67679;
  wire net_67680;
  wire net_67681;
  wire net_67684;
  wire net_67685;
  wire net_67686;
  wire net_67687;
  wire net_67691;
  wire net_67693;
  wire net_67696;
  wire net_67697;
  wire net_67698;
  wire net_67699;
  wire net_67702;
  wire net_67703;
  wire net_67704;
  wire net_67705;
  wire net_67708;
  wire net_67709;
  wire net_67710;
  wire net_67711;
  wire net_67712;
  wire net_67713;
  wire net_67720;
  wire net_67721;
  wire net_67722;
  wire net_67748;
  wire net_67757;
  wire net_67758;
  wire net_67759;
  wire net_67761;
  wire net_67765;
  wire net_67767;
  wire net_67770;
  wire net_67772;
  wire net_67774;
  wire net_67778;
  wire net_67789;
  wire net_67790;
  wire net_67791;
  wire net_67792;
  wire net_67802;
  wire net_67813;
  wire net_67814;
  wire net_67815;
  wire net_67816;
  wire net_67825;
  wire net_67827;
  wire net_67835;
  wire net_67836;
  wire net_67868;
  wire net_67961;
  wire net_68036;
  wire net_68042;
  wire net_68043;
  wire net_68044;
  wire net_68056;
  wire net_68058;
  wire net_68077;
  wire net_68093;
  wire net_68185;
  wire net_68599;
  wire net_68601;
  wire net_68638;
  wire net_68645;
  wire net_68646;
  wire net_68647;
  wire net_68648;
  wire net_68649;
  wire net_68650;
  wire net_68651;
  wire net_68655;
  wire net_68659;
  wire net_68662;
  wire net_68666;
  wire net_68670;
  wire net_68671;
  wire net_68675;
  wire net_68677;
  wire net_68680;
  wire net_68681;
  wire net_68687;
  wire net_68689;
  wire net_68698;
  wire net_68699;
  wire net_68701;
  wire net_68705;
  wire net_68706;
  wire net_68711;
  wire net_68712;
  wire net_68714;
  wire net_68715;
  wire net_68716;
  wire net_68717;
  wire net_68718;
  wire net_68719;
  wire net_68722;
  wire net_68723;
  wire net_68724;
  wire net_68758;
  wire net_68759;
  wire net_68764;
  wire net_68766;
  wire net_68768;
  wire net_68769;
  wire net_68771;
  wire net_68773;
  wire net_68774;
  wire net_68781;
  wire net_68782;
  wire net_68787;
  wire net_68792;
  wire net_68794;
  wire net_68815;
  wire net_68816;
  wire net_68817;
  wire net_68821;
  wire net_68822;
  wire net_68823;
  wire net_68824;
  wire net_68833;
  wire net_68834;
  wire net_68835;
  wire net_68836;
  wire net_68837;
  wire net_68838;
  wire net_68839;
  wire net_69120;
  wire net_69151;
  wire net_69166;
  wire net_69206;
  wire net_69207;
  wire net_69212;
  wire net_69347;
  wire net_69458;
  wire net_69461;
  wire net_69462;
  wire net_69503;
  wire net_69525;
  wire net_69535;
  wire net_69576;
  wire net_69577;
  wire net_69578;
  wire net_69579;
  wire net_69580;
  wire net_69581;
  wire net_69582;
  wire net_69583;
  wire net_69584;
  wire net_69585;
  wire net_69591;
  wire net_69606;
  wire net_69619;
  wire net_69623;
  wire net_69627;
  wire net_69629;
  wire net_69630;
  wire net_69670;
  wire net_69671;
  wire net_69673;
  wire net_69689;
  wire net_69690;
  wire net_69691;
  wire net_69698;
  wire net_69699;
  wire net_69700;
  wire net_69701;
  wire net_69702;
  wire net_69703;
  wire net_69704;
  wire net_69705;
  wire net_69706;
  wire net_69708;
  wire net_69713;
  wire net_69714;
  wire net_69716;
  wire net_69718;
  wire net_69722;
  wire net_69727;
  wire net_69742;
  wire net_69747;
  wire net_69749;
  wire net_69750;
  wire net_69753;
  wire net_69754;
  wire net_69756;
  wire net_69760;
  wire net_69763;
  wire net_69778;
  wire net_69788;
  wire net_69796;
  wire net_69802;
  wire net_69805;
  wire net_69806;
  wire net_69807;
  wire net_69808;
  wire net_69817;
  wire net_69822;
  wire net_69824;
  wire net_69826;
  wire net_69827;
  wire net_69828;
  wire net_69829;
  wire net_69830;
  wire net_69831;
  wire net_69847;
  wire net_69865;
  wire net_69867;
  wire net_69873;
  wire net_69875;
  wire net_69877;
  wire net_69878;
  wire net_69879;
  wire net_69880;
  wire net_69898;
  wire net_69900;
  wire net_69916;
  wire net_69918;
  wire net_69919;
  wire net_69923;
  wire net_69924;
  wire net_69925;
  wire net_69944;
  wire net_69945;
  wire net_69946;
  wire net_69949;
  wire net_69964;
  wire net_69967;
  wire net_69970;
  wire net_70003;
  wire net_70014;
  wire net_70017;
  wire net_70030;
  wire net_70065;
  wire net_70068;
  wire net_70069;
  wire net_70070;
  wire net_70071;
  wire net_70072;
  wire net_70073;
  wire net_70074;
  wire net_70075;
  wire net_70076;
  wire net_70077;
  wire net_70086;
  wire net_70093;
  wire net_70112;
  wire net_70113;
  wire net_70120;
  wire net_70121;
  wire net_70123;
  wire net_70124;
  wire net_70128;
  wire net_70136;
  wire net_70137;
  wire net_70138;
  wire net_70140;
  wire net_70145;
  wire net_70146;
  wire net_70147;
  wire net_70150;
  wire net_70151;
  wire net_70156;
  wire net_70157;
  wire net_70158;
  wire net_70175;
  wire net_70176;
  wire net_70186;
  wire net_70187;
  wire net_70188;
  wire net_70190;
  wire net_70191;
  wire net_70192;
  wire net_70195;
  wire net_70196;
  wire net_70197;
  wire net_70198;
  wire net_70199;
  wire net_70200;
  wire net_70206;
  wire net_70207;
  wire net_70209;
  wire net_70211;
  wire net_70236;
  wire net_70239;
  wire net_70243;
  wire net_70245;
  wire net_70247;
  wire net_70248;
  wire net_70254;
  wire net_70269;
  wire net_70274;
  wire net_70282;
  wire net_70288;
  wire net_70293;
  wire net_70305;
  wire net_70309;
  wire net_70314;
  wire net_70323;
  wire net_70324;
  wire net_70329;
  wire net_70344;
  wire net_70349;
  wire net_70350;
  wire net_70358;
  wire net_70362;
  wire net_70363;
  wire net_70365;
  wire net_70371;
  wire net_70374;
  wire net_70375;
  wire net_70376;
  wire net_70379;
  wire net_70382;
  wire net_70385;
  wire net_70388;
  wire net_70398;
  wire net_70414;
  wire net_70415;
  wire net_70416;
  wire net_70417;
  wire net_70420;
  wire net_70426;
  wire net_70427;
  wire net_70428;
  wire net_70429;
  wire net_70433;
  wire net_70434;
  wire net_70436;
  wire net_70437;
  wire net_70446;
  wire net_70461;
  wire net_70489;
  wire net_70493;
  wire net_70494;
  wire net_70497;
  wire net_70501;
  wire net_70502;
  wire net_70503;
  wire net_70507;
  wire net_70508;
  wire net_70515;
  wire net_70519;
  wire net_70520;
  wire net_70521;
  wire net_70522;
  wire net_70528;
  wire net_70543;
  wire net_70549;
  wire net_70550;
  wire net_70559;
  wire net_70560;
  wire net_70605;
  wire net_70606;
  wire net_70620;
  wire net_70668;
  wire net_70675;
  wire net_70682;
  wire net_70683;
  wire net_71574;
  wire net_71575;
  wire net_71577;
  wire net_71604;
  wire net_71608;
  wire net_71609;
  wire net_71614;
  wire net_71650;
  wire net_71651;
  wire net_71652;
  wire net_71653;
  wire net_71656;
  wire net_71657;
  wire net_71658;
  wire net_71659;
  wire net_71662;
  wire net_71663;
  wire net_71664;
  wire net_71665;
  wire net_71704;
  wire net_71794;
  wire net_71795;
  wire net_71837;
  wire net_71843;
  wire net_71844;
  wire net_71845;
  wire net_71851;
  wire net_71859;
  wire net_71867;
  wire net_71873;
  wire net_71874;
  wire net_71875;
  wire net_71878;
  wire net_71885;
  wire net_72466;
  wire net_72479;
  wire net_72484;
  wire net_72485;
  wire net_72495;
  wire net_72497;
  wire net_72530;
  wire net_72532;
  wire net_72541;
  wire net_72544;
  wire net_72545;
  wire net_72546;
  wire net_72547;
  wire net_72593;
  wire net_72594;
  wire net_72596;
  wire net_72597;
  wire net_72600;
  wire net_72601;
  wire net_72602;
  wire net_72604;
  wire net_72605;
  wire net_72607;
  wire net_72610;
  wire net_72612;
  wire net_72613;
  wire net_72618;
  wire net_72622;
  wire net_72624;
  wire net_72625;
  wire net_72628;
  wire net_72629;
  wire net_72630;
  wire net_72631;
  wire net_72635;
  wire net_72637;
  wire net_72652;
  wire net_72653;
  wire net_72654;
  wire net_72655;
  wire net_72659;
  wire net_72660;
  wire net_72661;
  wire net_72664;
  wire net_72666;
  wire net_72668;
  wire net_72669;
  wire net_72670;
  wire net_72685;
  wire net_72687;
  wire net_72692;
  wire net_73084;
  wire net_73085;
  wire net_73090;
  wire net_73105;
  wire net_73132;
  wire net_73133;
  wire net_73134;
  wire net_73135;
  wire net_73183;
  wire net_73330;
  wire net_73354;
  wire net_73355;
  wire net_73378;
  wire net_73396;
  wire net_73402;
  wire net_73407;
  wire net_73409;
  wire net_73410;
  wire net_73411;
  wire net_73412;
  wire net_73413;
  wire net_73414;
  wire net_73415;
  wire net_73416;
  wire net_73429;
  wire net_73439;
  wire net_73443;
  wire net_73452;
  wire net_73453;
  wire net_73454;
  wire net_73461;
  wire net_73462;
  wire net_73467;
  wire net_73473;
  wire net_73475;
  wire net_73478;
  wire net_73479;
  wire net_73481;
  wire net_73484;
  wire net_73492;
  wire net_73497;
  wire net_73502;
  wire net_73503;
  wire net_73504;
  wire net_73507;
  wire net_73509;
  wire net_73510;
  wire net_73514;
  wire net_73522;
  wire net_73527;
  wire net_73530;
  wire net_73532;
  wire net_73533;
  wire net_73534;
  wire net_73535;
  wire net_73536;
  wire net_73537;
  wire net_73538;
  wire net_73539;
  wire net_73544;
  wire net_73546;
  wire net_73550;
  wire net_73554;
  wire net_73560;
  wire net_73563;
  wire net_73574;
  wire net_73575;
  wire net_73576;
  wire net_73580;
  wire net_73582;
  wire net_73583;
  wire net_73585;
  wire net_73588;
  wire net_73589;
  wire net_73590;
  wire net_73591;
  wire net_73592;
  wire net_73595;
  wire net_73596;
  wire net_73599;
  wire net_73602;
  wire net_73604;
  wire net_73606;
  wire net_73607;
  wire net_73608;
  wire net_73613;
  wire net_73614;
  wire net_73615;
  wire net_73618;
  wire net_73619;
  wire net_73621;
  wire net_73624;
  wire net_73625;
  wire net_73627;
  wire net_73630;
  wire net_73632;
  wire net_73633;
  wire net_73636;
  wire net_73637;
  wire net_73639;
  wire net_73648;
  wire net_73650;
  wire net_73651;
  wire net_73652;
  wire net_73653;
  wire net_73654;
  wire net_73655;
  wire net_73656;
  wire net_73657;
  wire net_73658;
  wire net_73659;
  wire net_73660;
  wire net_73661;
  wire net_73662;
  wire net_73667;
  wire net_73669;
  wire net_73674;
  wire net_73675;
  wire net_73681;
  wire net_73701;
  wire net_73713;
  wire net_73717;
  wire net_73722;
  wire net_73723;
  wire net_73724;
  wire net_73725;
  wire net_73732;
  wire net_73744;
  wire net_73749;
  wire net_73753;
  wire net_73759;
  wire net_73767;
  wire net_73771;
  wire net_73776;
  wire net_73778;
  wire net_73779;
  wire net_73780;
  wire net_73781;
  wire net_73782;
  wire net_73783;
  wire net_73784;
  wire net_73785;
  wire net_73790;
  wire net_73795;
  wire net_73845;
  wire net_73849;
  wire net_73865;
  wire net_73867;
  wire net_73899;
  wire net_73901;
  wire net_73902;
  wire net_73903;
  wire net_73904;
  wire net_73905;
  wire net_73906;
  wire net_73907;
  wire net_73908;
  wire net_73919;
  wire net_73926;
  wire net_73946;
  wire net_73948;
  wire net_73950;
  wire net_73953;
  wire net_73955;
  wire net_73956;
  wire net_73962;
  wire net_73965;
  wire net_73969;
  wire net_73970;
  wire net_73971;
  wire net_73978;
  wire net_73983;
  wire net_73987;
  wire net_73994;
  wire net_74001;
  wire net_74005;
  wire net_74006;
  wire net_74007;
  wire net_74008;
  wire net_74013;
  wire net_74018;
  wire net_74022;
  wire net_74024;
  wire net_74025;
  wire net_74026;
  wire net_74027;
  wire net_74028;
  wire net_74029;
  wire net_74030;
  wire net_74031;
  wire net_74036;
  wire net_74038;
  wire net_74040;
  wire net_74042;
  wire net_74046;
  wire net_74047;
  wire net_74065;
  wire net_74068;
  wire net_74070;
  wire net_74072;
  wire net_74074;
  wire net_74076;
  wire net_74077;
  wire net_74080;
  wire net_74082;
  wire net_74083;
  wire net_74084;
  wire net_74086;
  wire net_74091;
  wire net_74092;
  wire net_74111;
  wire net_74112;
  wire net_74113;
  wire net_74116;
  wire net_74117;
  wire net_74119;
  wire net_74122;
  wire net_74124;
  wire net_74125;
  wire net_74128;
  wire net_74129;
  wire net_74131;
  wire net_74134;
  wire net_74135;
  wire net_74137;
  wire net_74140;
  wire net_74141;
  wire net_74143;
  wire net_74144;
  wire net_74145;
  wire net_74146;
  wire net_74165;
  wire net_74175;
  wire net_74195;
  wire net_74263;
  wire net_74267;
  wire net_74268;
  wire net_74300;
  wire net_74320;
  wire net_74387;
  wire net_74391;
  wire net_75655;
  wire net_75671;
  wire net_75674;
  wire net_75675;
  wire net_75676;
  wire net_75679;
  wire net_75682;
  wire net_76243;
  wire net_76245;
  wire net_76248;
  wire net_76250;
  wire net_76345;
  wire net_76391;
  wire net_76402;
  wire net_76408;
  wire net_76496;
  wire net_76508;
  wire net_76549;
  wire net_76550;
  wire net_76554;
  wire net_76651;
  wire net_76654;
  wire net_76656;
  wire net_76658;
  wire net_76699;
  wire net_76758;
  wire net_76795;
  wire net_76797;
  wire net_76800;
  wire net_76817;
  wire net_76855;
  wire net_76856;
  wire net_76857;
  wire net_76858;
  wire net_76859;
  wire net_76860;
  wire net_76861;
  wire net_76862;
  wire net_76911;
  wire net_76915;
  wire net_76919;
  wire net_76957;
  wire net_76958;
  wire net_76959;
  wire net_76960;
  wire net_76961;
  wire net_76962;
  wire net_76963;
  wire net_76964;
  wire net_77016;
  wire net_77027;
  wire net_77030;
  wire net_77031;
  wire net_77033;
  wire net_77034;
  wire net_77035;
  wire net_77036;
  wire net_77038;
  wire net_77039;
  wire net_77040;
  wire net_77042;
  wire net_77044;
  wire net_77048;
  wire net_77049;
  wire net_77050;
  wire net_77054;
  wire net_77056;
  wire net_77057;
  wire net_77059;
  wire net_77060;
  wire net_77061;
  wire net_77062;
  wire net_77063;
  wire net_77064;
  wire net_77065;
  wire net_77066;
  wire net_77075;
  wire net_77076;
  wire net_77078;
  wire net_77079;
  wire net_77080;
  wire net_77081;
  wire net_77082;
  wire net_77083;
  wire net_77086;
  wire net_77087;
  wire net_77088;
  wire net_77089;
  wire net_77090;
  wire net_77091;
  wire net_77092;
  wire net_77093;
  wire net_77094;
  wire net_77095;
  wire net_77096;
  wire net_77101;
  wire net_77110;
  wire net_77113;
  wire net_77114;
  wire net_77115;
  wire net_77116;
  wire net_77120;
  wire net_77122;
  wire net_77124;
  wire net_77129;
  wire net_77130;
  wire net_77131;
  wire net_77132;
  wire net_77133;
  wire net_77134;
  wire net_77135;
  wire net_77137;
  wire net_77141;
  wire net_77142;
  wire net_77147;
  wire net_77150;
  wire net_77151;
  wire net_77152;
  wire net_77156;
  wire net_77157;
  wire net_77158;
  wire net_77160;
  wire net_77161;
  wire net_77162;
  wire net_77163;
  wire net_77164;
  wire net_77165;
  wire net_77166;
  wire net_77167;
  wire net_77168;
  wire net_77177;
  wire net_77178;
  wire net_77180;
  wire net_77181;
  wire net_77182;
  wire net_77183;
  wire net_77184;
  wire net_77185;
  wire net_77188;
  wire net_77189;
  wire net_77190;
  wire net_77191;
  wire net_77192;
  wire net_77193;
  wire net_77194;
  wire net_77195;
  wire net_77196;
  wire net_77197;
  wire net_77198;
  wire net_77208;
  wire net_77217;
  wire net_77219;
  wire net_77220;
  wire net_77222;
  wire net_77223;
  wire net_77226;
  wire net_77231;
  wire net_77232;
  wire net_77233;
  wire net_77234;
  wire net_77235;
  wire net_77236;
  wire net_77239;
  wire net_77240;
  wire net_77246;
  wire net_77247;
  wire net_77248;
  wire net_77251;
  wire net_77252;
  wire net_77254;
  wire net_77258;
  wire net_77260;
  wire net_77261;
  wire net_77262;
  wire net_77264;
  wire net_77265;
  wire net_77266;
  wire net_77267;
  wire net_77268;
  wire net_77269;
  wire net_77270;
  wire net_77279;
  wire net_77280;
  wire net_77282;
  wire net_77283;
  wire net_77284;
  wire net_77285;
  wire net_77286;
  wire net_77287;
  wire net_77290;
  wire net_77291;
  wire net_77292;
  wire net_77293;
  wire net_77294;
  wire net_77295;
  wire net_77296;
  wire net_77297;
  wire net_77298;
  wire net_77299;
  wire net_77300;
  wire net_77322;
  wire net_77328;
  wire net_77334;
  wire net_77339;
  wire net_77342;
  wire net_77343;
  wire net_77346;
  wire net_77349;
  wire net_77351;
  wire net_77353;
  wire net_77354;
  wire net_77356;
  wire net_77357;
  wire net_77358;
  wire net_77359;
  wire net_77360;
  wire net_77361;
  wire net_77362;
  wire net_77363;
  wire net_77364;
  wire net_77365;
  wire net_77366;
  wire net_77367;
  wire net_77368;
  wire net_77369;
  wire net_77370;
  wire net_77371;
  wire net_77372;
  wire net_77381;
  wire net_77382;
  wire net_77384;
  wire net_77385;
  wire net_77386;
  wire net_77387;
  wire net_77388;
  wire net_77389;
  wire net_77392;
  wire net_77393;
  wire net_77394;
  wire net_77395;
  wire net_77396;
  wire net_77397;
  wire net_77398;
  wire net_77399;
  wire net_77400;
  wire net_77401;
  wire net_77402;
  wire net_77407;
  wire net_77421;
  wire net_77423;
  wire net_77435;
  wire net_77436;
  wire net_77437;
  wire net_77439;
  wire net_77440;
  wire net_77446;
  wire net_77447;
  wire net_77449;
  wire net_77450;
  wire net_77452;
  wire net_77453;
  wire net_77456;
  wire net_77457;
  wire net_77461;
  wire net_77462;
  wire net_77464;
  wire net_77466;
  wire net_77468;
  wire net_77470;
  wire net_77471;
  wire net_77472;
  wire net_77474;
  wire net_77483;
  wire net_77484;
  wire net_77486;
  wire net_77487;
  wire net_77488;
  wire net_77489;
  wire net_77490;
  wire net_77491;
  wire net_77494;
  wire net_77495;
  wire net_77496;
  wire net_77497;
  wire net_77498;
  wire net_77499;
  wire net_77500;
  wire net_77501;
  wire net_77503;
  wire net_77504;
  wire net_77509;
  wire net_77510;
  wire net_77512;
  wire net_77513;
  wire net_77514;
  wire net_77516;
  wire net_77518;
  wire net_77538;
  wire net_77539;
  wire net_77541;
  wire net_77542;
  wire net_77545;
  wire net_77548;
  wire net_77549;
  wire net_77550;
  wire net_77553;
  wire net_77555;
  wire net_77558;
  wire net_77559;
  wire net_77561;
  wire net_77562;
  wire net_77563;
  wire net_77564;
  wire net_77565;
  wire net_77568;
  wire net_77575;
  wire net_77576;
  wire net_77585;
  wire net_77586;
  wire net_77588;
  wire net_77589;
  wire net_77590;
  wire net_77591;
  wire net_77592;
  wire net_77593;
  wire net_77596;
  wire net_77597;
  wire net_77598;
  wire net_77599;
  wire net_77600;
  wire net_77601;
  wire net_77602;
  wire net_77603;
  wire net_77604;
  wire net_77605;
  wire net_77606;
  wire net_79368;
  wire net_79480;
  wire net_79582;
  wire net_79584;
  wire net_79589;
  wire net_79611;
  wire net_79622;
  wire net_79624;
  wire net_79628;
  wire net_79630;
  wire net_79635;
  wire net_79638;
  wire net_79641;
  wire net_79646;
  wire net_79649;
  wire net_79653;
  wire net_79654;
  wire net_79655;
  wire net_79656;
  wire net_79667;
  wire net_79668;
  wire net_79685;
  wire net_79686;
  wire net_79697;
  wire net_79699;
  wire net_79700;
  wire net_79701;
  wire net_79720;
  wire net_79732;
  wire net_79734;
  wire net_79756;
  wire net_79761;
  wire net_79776;
  wire net_79778;
  wire net_79856;
  wire net_79948;
  wire net_79950;
  wire net_79954;
  wire net_79975;
  wire net_79978;
  wire net_79980;
  wire net_79991;
  wire net_79997;
  wire net_80000;
  wire net_80004;
  wire net_80014;
  wire net_80022;
  wire net_80025;
  wire net_80028;
  wire net_80053;
  wire net_80055;
  wire net_80068;
  wire net_80069;
  wire net_80071;
  wire net_80072;
  wire net_80075;
  wire net_80076;
  wire net_80094;
  wire net_80095;
  wire net_80096;
  wire net_80101;
  wire net_80106;
  wire net_80114;
  wire net_80117;
  wire net_80119;
  wire net_80121;
  wire net_80122;
  wire net_80123;
  wire net_80125;
  wire net_80129;
  wire net_80132;
  wire net_80136;
  wire net_80137;
  wire net_80139;
  wire net_80140;
  wire net_80146;
  wire net_80147;
  wire net_80148;
  wire net_80163;
  wire net_80164;
  wire net_80165;
  wire net_80166;
  wire net_80175;
  wire net_80176;
  wire net_80177;
  wire net_80178;
  wire net_80187;
  wire net_80189;
  wire net_80191;
  wire net_80192;
  wire net_80193;
  wire net_80206;
  wire net_80208;
  wire net_80215;
  wire net_80222;
  wire net_80229;
  wire net_80242;
  wire net_80300;
  wire net_80315;
  wire net_80319;
  wire net_80322;
  wire net_80324;
  wire net_80359;
  wire net_80360;
  wire net_80364;
  wire net_80368;
  wire net_80369;
  wire net_80371;
  wire net_80372;
  wire net_80373;
  wire net_80375;
  wire net_80376;
  wire net_80377;
  wire net_80378;
  wire net_80379;
  wire net_80380;
  wire net_80381;
  wire net_80385;
  wire net_80388;
  wire net_80389;
  wire net_80392;
  wire net_80393;
  wire net_80394;
  wire net_80397;
  wire net_80398;
  wire net_80400;
  wire net_80404;
  wire net_80405;
  wire net_80406;
  wire net_80409;
  wire net_80410;
  wire net_80412;
  wire net_80415;
  wire net_80417;
  wire net_80418;
  wire net_80421;
  wire net_80422;
  wire net_80424;
  wire net_80428;
  wire net_80429;
  wire net_80430;
  wire net_80433;
  wire net_80435;
  wire net_80436;
  wire net_80437;
  wire net_80438;
  wire net_80439;
  wire net_80440;
  wire net_80441;
  wire net_80442;
  wire net_80443;
  wire net_80444;
  wire net_80446;
  wire net_80447;
  wire net_80464;
  wire net_80470;
  wire net_80473;
  wire net_80481;
  wire net_80482;
  wire net_80483;
  wire net_80485;
  wire net_80486;
  wire net_80489;
  wire net_80491;
  wire net_80492;
  wire net_80493;
  wire net_80494;
  wire net_80495;
  wire net_80499;
  wire net_80501;
  wire net_80502;
  wire net_80503;
  wire net_80507;
  wire net_80509;
  wire net_80510;
  wire net_80511;
  wire net_80514;
  wire net_80515;
  wire net_80516;
  wire net_80517;
  wire net_80521;
  wire net_80522;
  wire net_80523;
  wire net_80526;
  wire net_80528;
  wire net_80529;
  wire net_80532;
  wire net_80533;
  wire net_80535;
  wire net_80538;
  wire net_80539;
  wire net_80540;
  wire net_80544;
  wire net_80545;
  wire net_80547;
  wire net_80550;
  wire net_80551;
  wire net_80552;
  wire net_80556;
  wire net_80557;
  wire net_80558;
  wire net_80560;
  wire net_80561;
  wire net_80562;
  wire net_80563;
  wire net_80564;
  wire net_80565;
  wire net_80566;
  wire net_80567;
  wire net_80568;
  wire net_80569;
  wire net_80570;
  wire net_80589;
  wire net_80596;
  wire net_80604;
  wire net_80605;
  wire net_80609;
  wire net_80611;
  wire net_80612;
  wire net_80613;
  wire net_80618;
  wire net_80619;
  wire net_80620;
  wire net_80622;
  wire net_80623;
  wire net_80624;
  wire net_80626;
  wire net_80628;
  wire net_80631;
  wire net_80635;
  wire net_80637;
  wire net_80638;
  wire net_80639;
  wire net_80644;
  wire net_80649;
  wire net_80655;
  wire net_80656;
  wire net_80657;
  wire net_80658;
  wire net_80664;
  wire net_80667;
  wire net_80669;
  wire net_80670;
  wire net_80673;
  wire net_80674;
  wire net_80676;
  wire net_80679;
  wire net_80680;
  wire net_80681;
  wire net_80682;
  wire net_80684;
  wire net_80686;
  wire net_80687;
  wire net_80688;
  wire net_80689;
  wire net_80690;
  wire net_80691;
  wire net_80692;
  wire net_80693;
  wire net_80710;
  wire net_80718;
  wire net_80727;
  wire net_80729;
  wire net_80731;
  wire net_80735;
  wire net_80736;
  wire net_80738;
  wire net_80739;
  wire net_80740;
  wire net_80741;
  wire net_80743;
  wire net_80744;
  wire net_80745;
  wire net_80747;
  wire net_80749;
  wire net_80751;
  wire net_80752;
  wire net_80753;
  wire net_80755;
  wire net_80757;
  wire net_80760;
  wire net_80761;
  wire net_80762;
  wire net_80767;
  wire net_80768;
  wire net_80769;
  wire net_80772;
  wire net_80774;
  wire net_80775;
  wire net_80778;
  wire net_80779;
  wire net_80780;
  wire net_80784;
  wire net_80785;
  wire net_80787;
  wire net_80790;
  wire net_80791;
  wire net_80793;
  wire net_80797;
  wire net_80798;
  wire net_80799;
  wire net_80802;
  wire net_80804;
  wire net_80805;
  wire net_80806;
  wire net_80807;
  wire net_80808;
  wire net_80812;
  wire net_80813;
  wire net_80815;
  wire net_80833;
  wire net_80835;
  wire net_80838;
  wire net_80839;
  wire net_80844;
  wire net_80855;
  wire net_80859;
  wire net_80862;
  wire net_80864;
  wire net_80868;
  wire net_80870;
  wire net_80871;
  wire net_80877;
  wire net_80881;
  wire net_80882;
  wire net_80884;
  wire net_80885;
  wire net_80888;
  wire net_80890;
  wire net_80892;
  wire net_80894;
  wire net_80897;
  wire net_80898;
  wire net_80900;
  wire net_80902;
  wire net_80904;
  wire net_80906;
  wire net_80908;
  wire net_80910;
  wire net_80912;
  wire net_80915;
  wire net_80916;
  wire net_80918;
  wire net_80920;
  wire net_80922;
  wire net_80926;
  wire net_80928;
  wire net_80930;
  wire net_80932;
  wire net_80933;
  wire net_80934;
  wire net_80935;
  wire net_80936;
  wire net_80937;
  wire net_80938;
  wire net_80939;
  wire net_80950;
  wire net_80958;
  wire net_80963;
  wire net_80975;
  wire net_80976;
  wire net_80977;
  wire net_80978;
  wire net_80979;
  wire net_80980;
  wire net_80984;
  wire net_80985;
  wire net_80986;
  wire net_80987;
  wire net_80989;
  wire net_80990;
  wire net_80991;
  wire net_80992;
  wire net_80993;
  wire net_80995;
  wire net_80996;
  wire net_80997;
  wire net_80998;
  wire net_81001;
  wire net_81002;
  wire net_81003;
  wire net_81006;
  wire net_81007;
  wire net_81008;
  wire net_81009;
  wire net_81012;
  wire net_81014;
  wire net_81015;
  wire net_81018;
  wire net_81019;
  wire net_81020;
  wire net_81021;
  wire net_81024;
  wire net_81025;
  wire net_81027;
  wire net_81030;
  wire net_81031;
  wire net_81032;
  wire net_81033;
  wire net_81036;
  wire net_81038;
  wire net_81039;
  wire net_81043;
  wire net_81044;
  wire net_81045;
  wire net_81048;
  wire net_81050;
  wire net_81051;
  wire net_81052;
  wire net_81053;
  wire net_81054;
  wire net_81055;
  wire net_81056;
  wire net_81057;
  wire net_81058;
  wire net_81059;
  wire net_81060;
  wire net_81061;
  wire net_81062;
  wire net_81068;
  wire net_81081;
  wire net_81098;
  wire net_81099;
  wire net_81102;
  wire net_81103;
  wire net_81105;
  wire net_81107;
  wire net_81110;
  wire net_81111;
  wire net_81112;
  wire net_81115;
  wire net_81119;
  wire net_81120;
  wire net_81125;
  wire net_81135;
  wire net_81136;
  wire net_81138;
  wire net_81148;
  wire net_81149;
  wire net_81150;
  wire net_81153;
  wire net_81154;
  wire net_81155;
  wire net_81159;
  wire net_81160;
  wire net_81161;
  wire net_81162;
  wire net_81172;
  wire net_81173;
  wire net_81174;
  wire net_81175;
  wire net_81176;
  wire net_81177;
  wire net_81180;
  wire net_81181;
  wire net_81236;
  wire net_81240;
  wire net_81289;
  wire net_81294;
  wire net_81299;
  wire net_82776;
  wire net_83194;
  wire net_83198;
  wire net_83456;
  wire net_83460;
  wire net_83466;
  wire net_83503;
  wire net_83504;
  wire net_83505;
  wire net_83514;
  wire net_83515;
  wire net_83547;
  wire net_83564;
  wire net_83666;
  wire net_83667;
  wire net_83780;
  wire net_83822;
  wire net_83828;
  wire net_83833;
  wire net_83835;
  wire net_83843;
  wire net_83849;
  wire net_83854;
  wire net_83855;
  wire net_83866;
  wire net_83867;
  wire net_83889;
  wire net_83890;
  wire net_83892;
  wire net_83899;
  wire net_83900;
  wire net_83901;
  wire net_83914;
  wire net_83926;
  wire net_83943;
  wire net_83945;
  wire net_83946;
  wire net_83947;
  wire net_83956;
  wire net_83963;
  wire net_83964;
  wire net_83967;
  wire net_83972;
  wire net_83976;
  wire net_83978;
  wire net_83982;
  wire net_83985;
  wire net_84001;
  wire net_84002;
  wire net_84006;
  wire net_84007;
  wire net_84009;
  wire net_84022;
  wire net_84023;
  wire net_84024;
  wire net_84039;
  wire net_84041;
  wire net_84047;
  wire net_84189;
  wire net_84196;
  wire net_84197;
  wire net_84202;
  wire net_84204;
  wire net_84217;
  wire net_84235;
  wire net_84252;
  wire net_84253;
  wire net_84254;
  wire net_84255;
  wire net_84267;
  wire net_84269;
  wire net_84273;
  wire net_84276;
  wire net_84313;
  wire net_84314;
  wire net_84316;
  wire net_84319;
  wire net_84321;
  wire net_84322;
  wire net_84324;
  wire net_84325;
  wire net_84326;
  wire net_84327;
  wire net_84328;
  wire net_84333;
  wire net_84334;
  wire net_84335;
  wire net_84338;
  wire net_84341;
  wire net_84342;
  wire net_84343;
  wire net_84345;
  wire net_84346;
  wire net_84347;
  wire net_84351;
  wire net_84352;
  wire net_84353;
  wire net_84357;
  wire net_84358;
  wire net_84359;
  wire net_84360;
  wire net_84363;
  wire net_84364;
  wire net_84366;
  wire net_84369;
  wire net_84370;
  wire net_84371;
  wire net_84381;
  wire net_84382;
  wire net_84383;
  wire net_84387;
  wire net_84388;
  wire net_84390;
  wire net_84391;
  wire net_84392;
  wire net_84393;
  wire net_84397;
  wire net_84423;
  wire net_84436;
  wire net_84437;
  wire net_84438;
  wire net_84439;
  wire net_84441;
  wire net_84442;
  wire net_84443;
  wire net_84444;
  wire net_84445;
  wire net_84446;
  wire net_84447;
  wire net_84448;
  wire net_84450;
  wire net_84452;
  wire net_84453;
  wire net_84454;
  wire net_84455;
  wire net_84456;
  wire net_84458;
  wire net_84459;
  wire net_84462;
  wire net_84463;
  wire net_84465;
  wire net_84466;
  wire net_84468;
  wire net_84474;
  wire net_84475;
  wire net_84476;
  wire net_84477;
  wire net_84480;
  wire net_84481;
  wire net_84482;
  wire net_84483;
  wire net_84486;
  wire net_84487;
  wire net_84488;
  wire net_84489;
  wire net_84492;
  wire net_84493;
  wire net_84494;
  wire net_84495;
  wire net_84498;
  wire net_84499;
  wire net_84500;
  wire net_84501;
  wire net_84504;
  wire net_84505;
  wire net_84506;
  wire net_84507;
  wire net_84510;
  wire net_84511;
  wire net_84512;
  wire net_84513;
  wire net_84514;
  wire net_84515;
  wire net_84519;
  wire net_84521;
  wire net_84544;
  wire net_84548;
  wire net_84550;
  wire net_84558;
  wire net_84560;
  wire net_84561;
  wire net_84562;
  wire net_84563;
  wire net_84564;
  wire net_84566;
  wire net_84567;
  wire net_84568;
  wire net_84569;
  wire net_84570;
  wire net_84571;
  wire net_84572;
  wire net_84573;
  wire net_84575;
  wire net_84578;
  wire net_84581;
  wire net_84582;
  wire net_84583;
  wire net_84584;
  wire net_84585;
  wire net_84586;
  wire net_84589;
  wire net_84591;
  wire net_84592;
  wire net_84593;
  wire net_84594;
  wire net_84597;
  wire net_84598;
  wire net_84599;
  wire net_84600;
  wire net_84603;
  wire net_84604;
  wire net_84605;
  wire net_84609;
  wire net_84610;
  wire net_84612;
  wire net_84615;
  wire net_84617;
  wire net_84618;
  wire net_84621;
  wire net_84622;
  wire net_84623;
  wire net_84624;
  wire net_84627;
  wire net_84628;
  wire net_84629;
  wire net_84630;
  wire net_84633;
  wire net_84634;
  wire net_84635;
  wire net_84636;
  wire net_84637;
  wire net_84638;
  wire net_84639;
  wire net_84647;
  wire net_84664;
  wire net_84665;
  wire net_84666;
  wire net_84682;
  wire net_84686;
  wire net_84694;
  wire net_84696;
  wire net_84698;
  wire net_84706;
  wire net_84711;
  wire net_84732;
  wire net_84733;
  wire net_84734;
  wire net_84735;
  wire net_84739;
  wire net_84741;
  wire net_84750;
  wire net_84760;
  wire net_84761;
  wire net_84764;
  wire net_84765;
  wire net_84766;
  wire net_84767;
  wire net_84768;
  wire net_84769;
  wire net_84770;
  wire net_84792;
  wire net_84798;
  wire net_84806;
  wire net_84808;
  wire net_84812;
  wire net_84813;
  wire net_84814;
  wire net_84815;
  wire net_84817;
  wire net_84821;
  wire net_84822;
  wire net_84824;
  wire net_84825;
  wire net_84826;
  wire net_84827;
  wire net_84829;
  wire net_84830;
  wire net_84831;
  wire net_84832;
  wire net_84833;
  wire net_84834;
  wire net_84835;
  wire net_84837;
  wire net_84838;
  wire net_84839;
  wire net_84840;
  wire net_84843;
  wire net_84844;
  wire net_84845;
  wire net_84846;
  wire net_84849;
  wire net_84850;
  wire net_84851;
  wire net_84852;
  wire net_84858;
  wire net_84863;
  wire net_84870;
  wire net_84873;
  wire net_84874;
  wire net_84875;
  wire net_84876;
  wire net_84882;
  wire net_84884;
  wire net_84899;
  wire net_84901;
  wire net_84903;
  wire net_84907;
  wire net_84928;
  wire net_84929;
  wire net_84930;
  wire net_84931;
  wire net_84935;
  wire net_84936;
  wire net_84938;
  wire net_84939;
  wire net_84940;
  wire net_84941;
  wire net_84952;
  wire net_84953;
  wire net_84955;
  wire net_84957;
  wire net_84963;
  wire net_84966;
  wire net_84972;
  wire net_84973;
  wire net_84975;
  wire net_84980;
  wire net_84984;
  wire net_84985;
  wire net_84987;
  wire net_84990;
  wire net_84991;
  wire net_84992;
  wire net_84993;
  wire net_84996;
  wire net_84997;
  wire net_84999;
  wire net_85002;
  wire net_85003;
  wire net_85004;
  wire net_85005;
  wire net_85006;
  wire net_85007;
  wire net_85064;
  wire net_85098;
  wire net_85103;
  wire net_85129;
  wire net_85130;
  wire net_86563;
  wire net_86579;
  wire net_87513;
  wire net_87612;
  wire net_87617;
  wire net_87652;
  wire net_87655;
  wire net_87669;
  wire net_87692;
  wire net_87730;
  wire net_87731;
  wire net_87732;
  wire net_88152;
  wire net_88166;
  wire net_88190;
  wire net_88208;
  wire net_88223;
  wire net_88270;
  wire net_88278;
  wire net_88279;
  wire net_88318;
  wire net_88319;
  wire net_88320;
  wire net_88345;
  wire net_88346;
  wire net_88347;
  wire net_88374;
  wire net_88376;
  wire net_88382;
  wire net_88417;
  wire net_88419;
  wire net_88437;
  wire net_88449;
  wire net_88469;
  wire net_88496;
  wire net_88534;
  wire net_88539;
  wire net_88588;
  wire net_88590;
  wire net_88591;
  wire net_88592;
  wire net_88593;
  wire net_88636;
  wire net_88638;
  wire net_88639;
  wire net_88640;
  wire net_88642;
  wire net_88646;
  wire net_88647;
  wire net_88650;
  wire net_88656;
  wire net_88667;
  wire net_88669;
  wire net_88670;
  wire net_88673;
  wire net_88676;
  wire net_88677;
  wire net_88679;
  wire net_88681;
  wire net_88683;
  wire net_88685;
  wire net_88687;
  wire net_88689;
  wire net_88691;
  wire net_88693;
  wire net_88695;
  wire net_88697;
  wire net_88699;
  wire net_88701;
  wire net_88703;
  wire net_88705;
  wire net_88707;
  wire net_88712;
  wire net_88713;
  wire net_88739;
  wire net_91484;
  wire net_91491;
  wire net_91493;
  wire net_91495;
  wire net_91506;
  wire net_91516;
  wire net_91520;
  wire net_91522;
  wire net_91529;
  wire net_91530;
  wire net_91557;
  wire net_91558;
  wire net_91560;
  wire net_91561;
  wire net_91562;
  wire net_91563;
  wire dangling_wire_0;
  wire dangling_wire_1;
  wire dangling_wire_10;
  wire dangling_wire_11;
  wire dangling_wire_12;
  wire dangling_wire_13;
  wire dangling_wire_14;
  wire dangling_wire_15;
  wire dangling_wire_16;
  wire dangling_wire_17;
  wire dangling_wire_18;
  wire dangling_wire_19;
  wire dangling_wire_2;
  wire dangling_wire_20;
  wire dangling_wire_21;
  wire dangling_wire_22;
  wire dangling_wire_23;
  wire dangling_wire_24;
  wire dangling_wire_25;
  wire dangling_wire_26;
  wire dangling_wire_27;
  wire dangling_wire_28;
  wire dangling_wire_29;
  wire dangling_wire_3;
  wire dangling_wire_30;
  wire dangling_wire_31;
  wire dangling_wire_32;
  wire dangling_wire_33;
  wire dangling_wire_34;
  wire dangling_wire_35;
  wire dangling_wire_36;
  wire dangling_wire_37;
  wire dangling_wire_38;
  wire dangling_wire_39;
  wire dangling_wire_4;
  wire dangling_wire_40;
  wire dangling_wire_41;
  wire dangling_wire_42;
  wire dangling_wire_43;
  wire dangling_wire_44;
  wire dangling_wire_45;
  wire dangling_wire_46;
  wire dangling_wire_47;
  wire dangling_wire_48;
  wire dangling_wire_49;
  wire dangling_wire_5;
  wire dangling_wire_50;
  wire dangling_wire_51;
  wire dangling_wire_52;
  wire dangling_wire_53;
  wire dangling_wire_54;
  wire dangling_wire_55;
  wire dangling_wire_56;
  wire dangling_wire_57;
  wire dangling_wire_58;
  wire dangling_wire_59;
  wire dangling_wire_6;
  wire dangling_wire_60;
  wire dangling_wire_61;
  wire dangling_wire_62;
  wire dangling_wire_63;
  wire dangling_wire_64;
  wire dangling_wire_65;
  wire dangling_wire_66;
  wire dangling_wire_7;
  wire dangling_wire_8;
  wire dangling_wire_9;
  wire net_12210;
  wire net_12213_cascademuxed;
  wire net_12216;
  wire net_12222;
  wire net_12225_cascademuxed;
  wire net_12231_cascademuxed;
  wire net_12243_cascademuxed;
  wire net_12249_cascademuxed;
  wire net_13560_cascademuxed;
  wire net_16656;
  wire net_16659_cascademuxed;
  wire net_16662;
  wire net_16665_cascademuxed;
  wire net_16668;
  wire net_16689_cascademuxed;
  wire net_16695_cascademuxed;
  wire net_17271;
  wire net_17277;
  wire net_17280_cascademuxed;
  wire net_17283;
  wire net_17286_cascademuxed;
  wire net_17289;
  wire net_17292_cascademuxed;
  wire net_17295;
  wire net_17298_cascademuxed;
  wire net_17301;
  wire net_17304_cascademuxed;
  wire net_17388;
  wire net_17394;
  wire net_17397_cascademuxed;
  wire net_17400;
  wire net_17406;
  wire net_17412;
  wire net_17415_cascademuxed;
  wire net_17418;
  wire net_17421_cascademuxed;
  wire net_17424;
  wire net_17427_cascademuxed;
  wire net_17433_cascademuxed;
  wire net_17511;
  wire net_17514_cascademuxed;
  wire net_17517;
  wire net_17523;
  wire net_17526_cascademuxed;
  wire net_17529;
  wire net_17535;
  wire net_17541;
  wire net_17544_cascademuxed;
  wire net_20514_cascademuxed;
  wire net_20982_cascademuxed;
  wire net_21099_cascademuxed;
  wire net_21111_cascademuxed;
  wire net_21135_cascademuxed;
  wire net_21141_cascademuxed;
  wire net_21228_cascademuxed;
  wire net_21234_cascademuxed;
  wire net_21246_cascademuxed;
  wire net_21351_cascademuxed;
  wire net_23331_cascademuxed;
  wire net_25188_cascademuxed;
  wire net_29836_cascademuxed;
  wire net_31223_cascademuxed;
  wire net_31226;
  wire net_31253_cascademuxed;
  wire net_33830_cascademuxed;
  wire net_33842_cascademuxed;
  wire net_33848_cascademuxed;
  wire net_33854_cascademuxed;
  wire net_33860_cascademuxed;
  wire net_33866_cascademuxed;
  wire net_33971_cascademuxed;
  wire net_33977_cascademuxed;
  wire net_33983_cascademuxed;
  wire net_34811;
  wire net_34817;
  wire net_34820_cascademuxed;
  wire net_34823;
  wire net_34838_cascademuxed;
  wire net_34844_cascademuxed;
  wire net_34850_cascademuxed;
  wire net_34961_cascademuxed;
  wire net_35060_cascademuxed;
  wire net_35699_cascademuxed;
  wire net_36656;
  wire net_36662;
  wire net_36665_cascademuxed;
  wire net_36668;
  wire net_36671_cascademuxed;
  wire net_36689_cascademuxed;
  wire net_36695_cascademuxed;
  wire net_37655_cascademuxed;
  wire net_37661_cascademuxed;
  wire net_37667_cascademuxed;
  wire net_37673_cascademuxed;
  wire net_37679_cascademuxed;
  wire net_37691_cascademuxed;
  wire net_37778_cascademuxed;
  wire net_37784_cascademuxed;
  wire net_37790_cascademuxed;
  wire net_37796_cascademuxed;
  wire net_37802_cascademuxed;
  wire net_37808_cascademuxed;
  wire net_37814_cascademuxed;
  wire net_37820_cascademuxed;
  wire net_37901_cascademuxed;
  wire net_37931_cascademuxed;
  wire net_38393_cascademuxed;
  wire net_38396;
  wire net_38402;
  wire net_38405_cascademuxed;
  wire net_38408;
  wire net_38411_cascademuxed;
  wire net_38414;
  wire net_38417_cascademuxed;
  wire net_38420;
  wire net_38423_cascademuxed;
  wire net_38429_cascademuxed;
  wire net_38645_cascademuxed;
  wire net_38675_cascademuxed;
  wire net_38681_cascademuxed;
  wire net_38891_cascademuxed;
  wire net_39629_cascademuxed;
  wire net_40736_cascademuxed;
  wire net_40760_cascademuxed;
  wire net_40859_cascademuxed;
  wire net_40865_cascademuxed;
  wire net_40889_cascademuxed;
  wire net_40976_cascademuxed;
  wire net_41006_cascademuxed;
  wire net_41099_cascademuxed;
  wire net_41111_cascademuxed;
  wire net_41489;
  wire net_41495;
  wire net_41501;
  wire net_41504_cascademuxed;
  wire net_41522_cascademuxed;
  wire net_41621_cascademuxed;
  wire net_41633_cascademuxed;
  wire net_41645_cascademuxed;
  wire net_41651_cascademuxed;
  wire net_42224_cascademuxed;
  wire net_42230_cascademuxed;
  wire net_42242_cascademuxed;
  wire net_42266_cascademuxed;
  wire net_42482_cascademuxed;
  wire net_42593_cascademuxed;
  wire net_42605_cascademuxed;
  wire net_42713;
  wire net_42716_cascademuxed;
  wire net_42719;
  wire net_42722_cascademuxed;
  wire net_42725;
  wire net_42728_cascademuxed;
  wire net_42731;
  wire net_42734_cascademuxed;
  wire net_42737;
  wire net_42740_cascademuxed;
  wire net_42743;
  wire net_42746_cascademuxed;
  wire net_42749;
  wire net_42752_cascademuxed;
  wire net_42758_cascademuxed;
  wire net_42836;
  wire net_42839_cascademuxed;
  wire net_42842;
  wire net_42845_cascademuxed;
  wire net_42848;
  wire net_42851_cascademuxed;
  wire net_42854;
  wire net_42857_cascademuxed;
  wire net_42860;
  wire net_42863_cascademuxed;
  wire net_42866;
  wire net_42869_cascademuxed;
  wire net_42875_cascademuxed;
  wire net_42881_cascademuxed;
  wire net_42962_cascademuxed;
  wire net_42974_cascademuxed;
  wire net_42992_cascademuxed;
  wire net_42998_cascademuxed;
  wire net_43085_cascademuxed;
  wire net_43109_cascademuxed;
  wire net_43331_cascademuxed;
  wire net_43334;
  wire net_43340;
  wire net_43346;
  wire net_43349_cascademuxed;
  wire net_43352;
  wire net_43355_cascademuxed;
  wire net_43358;
  wire net_43364;
  wire net_43367_cascademuxed;
  wire net_43451;
  wire net_43457;
  wire net_43460_cascademuxed;
  wire net_43463;
  wire net_43466_cascademuxed;
  wire net_43469;
  wire net_43475;
  wire net_43481;
  wire net_43484_cascademuxed;
  wire net_43487;
  wire net_43490_cascademuxed;
  wire net_43574;
  wire net_43580;
  wire net_43586;
  wire net_43589_cascademuxed;
  wire net_43592;
  wire net_43598;
  wire net_43604;
  wire net_43610;
  wire net_43613_cascademuxed;
  wire net_43619_cascademuxed;
  wire net_43697;
  wire net_43703;
  wire net_43706_cascademuxed;
  wire net_43718_cascademuxed;
  wire net_44561_cascademuxed;
  wire net_44564;
  wire net_44567_cascademuxed;
  wire net_44570;
  wire net_44576;
  wire net_44579_cascademuxed;
  wire net_44696_cascademuxed;
  wire net_44702_cascademuxed;
  wire net_44714_cascademuxed;
  wire net_44726_cascademuxed;
  wire net_44807_cascademuxed;
  wire net_44825_cascademuxed;
  wire net_44837_cascademuxed;
  wire net_44843_cascademuxed;
  wire net_44849_cascademuxed;
  wire net_44930_cascademuxed;
  wire net_44942_cascademuxed;
  wire net_44948_cascademuxed;
  wire net_44954_cascademuxed;
  wire net_44966_cascademuxed;
  wire net_44972_cascademuxed;
  wire net_45932_cascademuxed;
  wire net_45974_cascademuxed;
  wire net_46058;
  wire net_46061_cascademuxed;
  wire net_46064;
  wire net_46067_cascademuxed;
  wire net_46070;
  wire net_46073_cascademuxed;
  wire net_46076;
  wire net_46079_cascademuxed;
  wire net_46082;
  wire net_46085_cascademuxed;
  wire net_46091_cascademuxed;
  wire net_46097_cascademuxed;
  wire net_46202_cascademuxed;
  wire net_46208_cascademuxed;
  wire net_46214_cascademuxed;
  wire net_46220_cascademuxed;
  wire net_46301_cascademuxed;
  wire net_46319_cascademuxed;
  wire net_46331_cascademuxed;
  wire net_46337_cascademuxed;
  wire net_46436_cascademuxed;
  wire net_46553_cascademuxed;
  wire net_46565_cascademuxed;
  wire net_46571_cascademuxed;
  wire net_46670_cascademuxed;
  wire net_46676_cascademuxed;
  wire net_46682_cascademuxed;
  wire net_46688_cascademuxed;
  wire net_46694_cascademuxed;
  wire net_46700_cascademuxed;
  wire net_46706_cascademuxed;
  wire net_46712_cascademuxed;
  wire net_46805_cascademuxed;
  wire net_46823_cascademuxed;
  wire net_46829_cascademuxed;
  wire net_46835_cascademuxed;
  wire net_46940_cascademuxed;
  wire net_47069_cascademuxed;
  wire net_47168_cascademuxed;
  wire net_47291_cascademuxed;
  wire net_47297_cascademuxed;
  wire net_47420_cascademuxed;
  wire net_47543_cascademuxed;
  wire net_47936_cascademuxed;
  wire net_48668_cascademuxed;
  wire net_48767_cascademuxed;
  wire net_48779_cascademuxed;
  wire net_49892_cascademuxed;
  wire net_49922_cascademuxed;
  wire net_50261_cascademuxed;
  wire net_50273_cascademuxed;
  wire net_50375;
  wire net_50378_cascademuxed;
  wire net_50381;
  wire net_50384_cascademuxed;
  wire net_50387;
  wire net_50390_cascademuxed;
  wire net_50393;
  wire net_50396_cascademuxed;
  wire net_50399;
  wire net_50402_cascademuxed;
  wire net_50405;
  wire net_50408_cascademuxed;
  wire net_50411;
  wire net_50414_cascademuxed;
  wire net_50420_cascademuxed;
  wire net_50498;
  wire net_50501_cascademuxed;
  wire net_50504;
  wire net_50507_cascademuxed;
  wire net_50510;
  wire net_50513_cascademuxed;
  wire net_50516;
  wire net_50519_cascademuxed;
  wire net_50522;
  wire net_50525_cascademuxed;
  wire net_50528;
  wire net_50531_cascademuxed;
  wire net_50537_cascademuxed;
  wire net_50543_cascademuxed;
  wire net_50624_cascademuxed;
  wire net_50636_cascademuxed;
  wire net_50654_cascademuxed;
  wire net_50666_cascademuxed;
  wire net_50759_cascademuxed;
  wire net_50771_cascademuxed;
  wire net_50777_cascademuxed;
  wire net_50789_cascademuxed;
  wire net_50876_cascademuxed;
  wire net_50906_cascademuxed;
  wire net_50993_cascademuxed;
  wire net_50999_cascademuxed;
  wire net_51116_cascademuxed;
  wire net_51128_cascademuxed;
  wire net_51251_cascademuxed;
  wire net_51263_cascademuxed;
  wire net_51485_cascademuxed;
  wire net_51521_cascademuxed;
  wire net_51527_cascademuxed;
  wire net_52223_cascademuxed;
  wire net_52226;
  wire net_52229_cascademuxed;
  wire net_52232;
  wire net_52238;
  wire net_52241_cascademuxed;
  wire net_52352_cascademuxed;
  wire net_52358_cascademuxed;
  wire net_53144_cascademuxed;
  wire net_53225_cascademuxed;
  wire net_53228;
  wire net_53231_cascademuxed;
  wire net_53234;
  wire net_53237_cascademuxed;
  wire net_53240;
  wire net_53255_cascademuxed;
  wire net_53267_cascademuxed;
  wire net_53720;
  wire net_53726;
  wire net_53732;
  wire net_53735_cascademuxed;
  wire net_53738;
  wire net_53741_cascademuxed;
  wire net_53744;
  wire net_53747_cascademuxed;
  wire net_53753_cascademuxed;
  wire net_53759_cascademuxed;
  wire net_53840_cascademuxed;
  wire net_53846_cascademuxed;
  wire net_53852_cascademuxed;
  wire net_53870_cascademuxed;
  wire net_53876_cascademuxed;
  wire net_54209_cascademuxed;
  wire net_54215_cascademuxed;
  wire net_54221_cascademuxed;
  wire net_54227_cascademuxed;
  wire net_54245_cascademuxed;
  wire net_54332_cascademuxed;
  wire net_54338_cascademuxed;
  wire net_54344_cascademuxed;
  wire net_54356_cascademuxed;
  wire net_54374_cascademuxed;
  wire net_54455_cascademuxed;
  wire net_54461_cascademuxed;
  wire net_54467_cascademuxed;
  wire net_54473_cascademuxed;
  wire net_54491_cascademuxed;
  wire net_54578_cascademuxed;
  wire net_54596_cascademuxed;
  wire net_54614_cascademuxed;
  wire net_54620_cascademuxed;
  wire net_54698;
  wire net_54701_cascademuxed;
  wire net_54704;
  wire net_54707_cascademuxed;
  wire net_54710;
  wire net_54713_cascademuxed;
  wire net_54716;
  wire net_54719_cascademuxed;
  wire net_54722;
  wire net_54725_cascademuxed;
  wire net_54728;
  wire net_54731_cascademuxed;
  wire net_54734;
  wire net_54737_cascademuxed;
  wire net_54743_cascademuxed;
  wire net_54821;
  wire net_54824_cascademuxed;
  wire net_54827;
  wire net_54830_cascademuxed;
  wire net_54833;
  wire net_54836_cascademuxed;
  wire net_54839;
  wire net_54842_cascademuxed;
  wire net_54845;
  wire net_54848_cascademuxed;
  wire net_54851;
  wire net_54854_cascademuxed;
  wire net_54860_cascademuxed;
  wire net_54866_cascademuxed;
  wire net_55076_cascademuxed;
  wire net_55082_cascademuxed;
  wire net_55094_cascademuxed;
  wire net_55106_cascademuxed;
  wire net_55112_cascademuxed;
  wire net_55217_cascademuxed;
  wire net_55223_cascademuxed;
  wire net_55229_cascademuxed;
  wire net_55235_cascademuxed;
  wire net_55457_cascademuxed;
  wire net_55481_cascademuxed;
  wire net_56066_cascademuxed;
  wire net_56084_cascademuxed;
  wire net_56090_cascademuxed;
  wire net_56821_cascademuxed;
  wire net_56827_cascademuxed;
  wire net_56839_cascademuxed;
  wire net_56845_cascademuxed;
  wire net_56932_cascademuxed;
  wire net_56938_cascademuxed;
  wire net_56950_cascademuxed;
  wire net_56956_cascademuxed;
  wire net_56962_cascademuxed;
  wire net_56968_cascademuxed;
  wire net_57061_cascademuxed;
  wire net_57085_cascademuxed;
  wire net_57097_cascademuxed;
  wire net_57430_cascademuxed;
  wire net_57460_cascademuxed;
  wire net_57466_cascademuxed;
  wire net_57571_cascademuxed;
  wire net_57583_cascademuxed;
  wire net_57589_cascademuxed;
  wire net_57673;
  wire net_57676_cascademuxed;
  wire net_57679;
  wire net_57682_cascademuxed;
  wire net_57685;
  wire net_57688_cascademuxed;
  wire net_57691;
  wire net_57694_cascademuxed;
  wire net_57697;
  wire net_57700_cascademuxed;
  wire net_57706_cascademuxed;
  wire net_57712_cascademuxed;
  wire net_57835_cascademuxed;
  wire net_57928_cascademuxed;
  wire net_57940_cascademuxed;
  wire net_57952_cascademuxed;
  wire net_58039_cascademuxed;
  wire net_58051_cascademuxed;
  wire net_58057_cascademuxed;
  wire net_58081_cascademuxed;
  wire net_58168_cascademuxed;
  wire net_58174_cascademuxed;
  wire net_58180_cascademuxed;
  wire net_58186_cascademuxed;
  wire net_58192_cascademuxed;
  wire net_58198_cascademuxed;
  wire net_58285_cascademuxed;
  wire net_58291_cascademuxed;
  wire net_58297_cascademuxed;
  wire net_58309_cascademuxed;
  wire net_58315_cascademuxed;
  wire net_58327_cascademuxed;
  wire net_58414_cascademuxed;
  wire net_58420_cascademuxed;
  wire net_58426_cascademuxed;
  wire net_58432_cascademuxed;
  wire net_58438_cascademuxed;
  wire net_58531_cascademuxed;
  wire net_58537_cascademuxed;
  wire net_58555_cascademuxed;
  wire net_58801_cascademuxed;
  wire net_58819_cascademuxed;
  wire net_58906_cascademuxed;
  wire net_58936_cascademuxed;
  wire net_59023_cascademuxed;
  wire net_59029_cascademuxed;
  wire net_59035_cascademuxed;
  wire net_59053_cascademuxed;
  wire net_59065_cascademuxed;
  wire net_59785_cascademuxed;
  wire net_59890_cascademuxed;
  wire net_59914_cascademuxed;
  wire net_60639_cascademuxed;
  wire net_60645_cascademuxed;
  wire net_60651_cascademuxed;
  wire net_60657_cascademuxed;
  wire net_60768_cascademuxed;
  wire net_60786_cascademuxed;
  wire net_60792_cascademuxed;
  wire net_60798_cascademuxed;
  wire net_60804_cascademuxed;
  wire net_61530_cascademuxed;
  wire net_61542_cascademuxed;
  wire net_61623_cascademuxed;
  wire net_61629_cascademuxed;
  wire net_61647_cascademuxed;
  wire net_61653_cascademuxed;
  wire net_61659_cascademuxed;
  wire net_61743;
  wire net_61746_cascademuxed;
  wire net_61749;
  wire net_61752_cascademuxed;
  wire net_61755;
  wire net_61758_cascademuxed;
  wire net_61761;
  wire net_61764_cascademuxed;
  wire net_61767;
  wire net_61770_cascademuxed;
  wire net_61773;
  wire net_61776_cascademuxed;
  wire net_61779;
  wire net_61782_cascademuxed;
  wire net_61788_cascademuxed;
  wire net_61866;
  wire net_61869_cascademuxed;
  wire net_61872;
  wire net_61875_cascademuxed;
  wire net_61878;
  wire net_61881_cascademuxed;
  wire net_61884;
  wire net_61887_cascademuxed;
  wire net_61890;
  wire net_61893_cascademuxed;
  wire net_61896;
  wire net_61899_cascademuxed;
  wire net_61905_cascademuxed;
  wire net_61911_cascademuxed;
  wire net_61992_cascademuxed;
  wire net_61998_cascademuxed;
  wire net_62004_cascademuxed;
  wire net_62010_cascademuxed;
  wire net_62022_cascademuxed;
  wire net_62028_cascademuxed;
  wire net_62034_cascademuxed;
  wire net_62121_cascademuxed;
  wire net_62139_cascademuxed;
  wire net_62145_cascademuxed;
  wire net_62157_cascademuxed;
  wire net_62250_cascademuxed;
  wire net_62256_cascademuxed;
  wire net_62262_cascademuxed;
  wire net_62268_cascademuxed;
  wire net_62280_cascademuxed;
  wire net_62385_cascademuxed;
  wire net_62403_cascademuxed;
  wire net_62484_cascademuxed;
  wire net_62490_cascademuxed;
  wire net_62502_cascademuxed;
  wire net_62526_cascademuxed;
  wire net_62607_cascademuxed;
  wire net_62613_cascademuxed;
  wire net_62619_cascademuxed;
  wire net_62643_cascademuxed;
  wire net_62748_cascademuxed;
  wire net_62766_cascademuxed;
  wire net_62865_cascademuxed;
  wire net_62889_cascademuxed;
  wire net_62895_cascademuxed;
  wire net_63228_cascademuxed;
  wire net_63252_cascademuxed;
  wire net_63264_cascademuxed;
  wire net_63837_cascademuxed;
  wire net_63861_cascademuxed;
  wire net_63867_cascademuxed;
  wire net_63879_cascademuxed;
  wire net_63990_cascademuxed;
  wire net_64002_cascademuxed;
  wire net_64488_cascademuxed;
  wire net_64500_cascademuxed;
  wire net_64842;
  wire net_64845_cascademuxed;
  wire net_64848;
  wire net_64854;
  wire net_64860;
  wire net_64866;
  wire net_64872;
  wire net_64962_cascademuxed;
  wire net_65343_cascademuxed;
  wire net_65355_cascademuxed;
  wire net_65361_cascademuxed;
  wire net_65367_cascademuxed;
  wire net_65583_cascademuxed;
  wire net_65700_cascademuxed;
  wire net_65706_cascademuxed;
  wire net_65712_cascademuxed;
  wire net_65730_cascademuxed;
  wire net_65736_cascademuxed;
  wire net_65835_cascademuxed;
  wire net_65952_cascademuxed;
  wire net_65976_cascademuxed;
  wire net_66069_cascademuxed;
  wire net_66081_cascademuxed;
  wire net_66087_cascademuxed;
  wire net_66099_cascademuxed;
  wire net_66105_cascademuxed;
  wire net_66198_cascademuxed;
  wire net_66321_cascademuxed;
  wire net_66450_cascademuxed;
  wire net_66456_cascademuxed;
  wire net_66567_cascademuxed;
  wire net_66585_cascademuxed;
  wire net_66591_cascademuxed;
  wire net_66597_cascademuxed;
  wire net_66690_cascademuxed;
  wire net_66696_cascademuxed;
  wire net_66702_cascademuxed;
  wire net_66708_cascademuxed;
  wire net_66714_cascademuxed;
  wire net_67674_cascademuxed;
  wire net_67680_cascademuxed;
  wire net_67686_cascademuxed;
  wire net_67698_cascademuxed;
  wire net_67704_cascademuxed;
  wire net_67710_cascademuxed;
  wire net_67791_cascademuxed;
  wire net_67815_cascademuxed;
  wire net_67827_cascademuxed;
  wire net_68670_cascademuxed;
  wire net_68706_cascademuxed;
  wire net_68712_cascademuxed;
  wire net_68817_cascademuxed;
  wire net_68823_cascademuxed;
  wire net_68835_cascademuxed;
  wire net_69690_cascademuxed;
  wire net_69807_cascademuxed;
  wire net_69900_cascademuxed;
  wire net_69918_cascademuxed;
  wire net_69924_cascademuxed;
  wire net_70065_cascademuxed;
  wire net_70146_cascademuxed;
  wire net_70158_cascademuxed;
  wire net_70176_cascademuxed;
  wire net_70188_cascademuxed;
  wire net_70269_cascademuxed;
  wire net_70293_cascademuxed;
  wire net_70305_cascademuxed;
  wire net_70398_cascademuxed;
  wire net_70416_cascademuxed;
  wire net_70428_cascademuxed;
  wire net_70434_cascademuxed;
  wire net_70515_cascademuxed;
  wire net_70521_cascademuxed;
  wire net_70668_cascademuxed;
  wire net_71652_cascademuxed;
  wire net_71658_cascademuxed;
  wire net_71664_cascademuxed;
  wire net_72624_cascademuxed;
  wire net_72630_cascademuxed;
  wire net_72654_cascademuxed;
  wire net_72660_cascademuxed;
  wire net_72666_cascademuxed;
  wire net_73134_cascademuxed;
  wire net_73497_cascademuxed;
  wire net_73503_cascademuxed;
  wire net_73509_cascademuxed;
  wire net_73527_cascademuxed;
  wire net_73608_cascademuxed;
  wire net_73614_cascademuxed;
  wire net_73632_cascademuxed;
  wire net_73650_cascademuxed;
  wire net_73749_cascademuxed;
  wire net_73767_cascademuxed;
  wire net_73983_cascademuxed;
  wire net_74001_cascademuxed;
  wire net_74007_cascademuxed;
  wire net_74013_cascademuxed;
  wire net_74112_cascademuxed;
  wire net_74124_cascademuxed;
  wire net_77075_cascademuxed;
  wire net_77076_cascademuxed;
  wire net_77078_cascademuxed;
  wire net_77079_cascademuxed;
  wire net_77080_cascademuxed;
  wire net_77081_cascademuxed;
  wire net_77082_cascademuxed;
  wire net_77083_cascademuxed;
  wire net_77177_cascademuxed;
  wire net_77178_cascademuxed;
  wire net_77180_cascademuxed;
  wire net_77181_cascademuxed;
  wire net_77182_cascademuxed;
  wire net_77183_cascademuxed;
  wire net_77184_cascademuxed;
  wire net_77185_cascademuxed;
  wire net_77279_cascademuxed;
  wire net_77280_cascademuxed;
  wire net_77282_cascademuxed;
  wire net_77283_cascademuxed;
  wire net_77284_cascademuxed;
  wire net_77285_cascademuxed;
  wire net_77286_cascademuxed;
  wire net_77287_cascademuxed;
  wire net_77381_cascademuxed;
  wire net_77382_cascademuxed;
  wire net_77384_cascademuxed;
  wire net_77385_cascademuxed;
  wire net_77386_cascademuxed;
  wire net_77387_cascademuxed;
  wire net_77388_cascademuxed;
  wire net_77389_cascademuxed;
  wire net_77483_cascademuxed;
  wire net_77484_cascademuxed;
  wire net_77486_cascademuxed;
  wire net_77487_cascademuxed;
  wire net_77488_cascademuxed;
  wire net_77489_cascademuxed;
  wire net_77490_cascademuxed;
  wire net_77491_cascademuxed;
  wire net_77585_cascademuxed;
  wire net_77586_cascademuxed;
  wire net_77588_cascademuxed;
  wire net_77589_cascademuxed;
  wire net_77590_cascademuxed;
  wire net_77591_cascademuxed;
  wire net_77592_cascademuxed;
  wire net_77593_cascademuxed;
  wire net_79655_cascademuxed;
  wire net_79667_cascademuxed;
  wire net_79685_cascademuxed;
  wire net_79697_cascademuxed;
  wire net_79778_cascademuxed;
  wire net_80147_cascademuxed;
  wire net_80165_cascademuxed;
  wire net_80177_cascademuxed;
  wire net_80189_cascademuxed;
  wire net_80300_cascademuxed;
  wire net_80393_cascademuxed;
  wire net_80405_cascademuxed;
  wire net_80417_cascademuxed;
  wire net_80429_cascademuxed;
  wire net_80435_cascademuxed;
  wire net_80516_cascademuxed;
  wire net_80522_cascademuxed;
  wire net_80528_cascademuxed;
  wire net_80540_cascademuxed;
  wire net_80552_cascademuxed;
  wire net_80558_cascademuxed;
  wire net_80639_cascademuxed;
  wire net_80657_cascademuxed;
  wire net_80669_cascademuxed;
  wire net_80681_cascademuxed;
  wire net_80762_cascademuxed;
  wire net_80768_cascademuxed;
  wire net_80774_cascademuxed;
  wire net_80780_cascademuxed;
  wire net_80798_cascademuxed;
  wire net_80804_cascademuxed;
  wire net_80882;
  wire net_80885_cascademuxed;
  wire net_80888;
  wire net_80894;
  wire net_80897_cascademuxed;
  wire net_80900;
  wire net_80906;
  wire net_80912;
  wire net_80915_cascademuxed;
  wire net_81008_cascademuxed;
  wire net_81014_cascademuxed;
  wire net_81020_cascademuxed;
  wire net_81032_cascademuxed;
  wire net_81038_cascademuxed;
  wire net_81044_cascademuxed;
  wire net_81050_cascademuxed;
  wire net_81149_cascademuxed;
  wire net_81155_cascademuxed;
  wire net_81161_cascademuxed;
  wire net_81173_cascademuxed;
  wire net_83504_cascademuxed;
  wire net_83855_cascademuxed;
  wire net_83867_cascademuxed;
  wire net_83978_cascademuxed;
  wire net_84002_cascademuxed;
  wire net_84254_cascademuxed;
  wire net_84347_cascademuxed;
  wire net_84353_cascademuxed;
  wire net_84359_cascademuxed;
  wire net_84371_cascademuxed;
  wire net_84383_cascademuxed;
  wire net_84476_cascademuxed;
  wire net_84482_cascademuxed;
  wire net_84488_cascademuxed;
  wire net_84494_cascademuxed;
  wire net_84500_cascademuxed;
  wire net_84506_cascademuxed;
  wire net_84512_cascademuxed;
  wire net_84593_cascademuxed;
  wire net_84599_cascademuxed;
  wire net_84605_cascademuxed;
  wire net_84617_cascademuxed;
  wire net_84623_cascademuxed;
  wire net_84629_cascademuxed;
  wire net_84635_cascademuxed;
  wire net_84734_cascademuxed;
  wire net_84839_cascademuxed;
  wire net_84845_cascademuxed;
  wire net_84851_cascademuxed;
  wire net_84863_cascademuxed;
  wire net_84875_cascademuxed;
  wire net_84980_cascademuxed;
  wire net_84992_cascademuxed;
  wire net_85004_cascademuxed;
  wire net_85103_cascademuxed;
  wire net_87692_cascademuxed;
  wire net_88190_cascademuxed;
  wire net_88208_cascademuxed;
  wire net_88319_cascademuxed;
  wire net_88667;
  wire net_88670_cascademuxed;
  wire net_88673;
  wire net_88676_cascademuxed;
  wire net_88679;
  wire net_88685;
  wire net_88691;
  wire net_88697;
  wire net_88712_cascademuxed;
  wire net_91529_cascademuxed;
  wire seg_10_10_local_g0_1_42436;
  wire seg_10_10_local_g0_6_42441;
  wire seg_10_10_lutff_2_out_38565;
  wire seg_10_10_neigh_op_lft_1_34733;
  wire seg_10_10_sp4_h_l_43_27633;
  wire seg_10_10_sp4_h_r_36_31037;
  wire seg_10_10_sp4_h_r_4_42535;
  wire seg_10_10_sp4_v_b_6_38348;
  wire seg_10_11_glb_netwk_0_5;
  wire seg_10_11_local_g0_2_42560;
  wire seg_10_11_local_g0_5_42563;
  wire seg_10_11_local_g2_2_42576;
  wire seg_10_11_local_g2_4_42578;
  wire seg_10_11_local_g2_7_42581;
  wire seg_10_11_local_g3_4_42586;
  wire seg_10_11_local_g3_5_42587;
  wire seg_10_11_lutff_0_out_38686;
  wire seg_10_11_lutff_1_out_38687;
  wire seg_10_11_lutff_4_out_38690;
  wire seg_10_11_neigh_op_bnl_4_34736;
  wire seg_10_11_neigh_op_bot_2_38565;
  wire seg_10_11_neigh_op_lft_5_34860;
  wire seg_10_11_neigh_op_rgt_2_42519;
  wire seg_10_11_neigh_op_rgt_7_42524;
  wire seg_10_11_sp4_r_v_b_21_42427;
  wire seg_10_11_sp4_r_v_b_37_42665;
  wire seg_10_12_glb_netwk_0_5;
  wire seg_10_12_local_g0_0_42681;
  wire seg_10_12_local_g0_1_42682;
  wire seg_10_12_local_g0_3_42684;
  wire seg_10_12_local_g0_4_42685;
  wire seg_10_12_local_g0_5_42686;
  wire seg_10_12_local_g0_6_42687;
  wire seg_10_12_local_g1_0_42689;
  wire seg_10_12_local_g1_1_42690;
  wire seg_10_12_local_g1_3_42692;
  wire seg_10_12_local_g1_4_42693;
  wire seg_10_12_local_g1_7_42696;
  wire seg_10_12_local_g2_1_42698;
  wire seg_10_12_local_g2_2_42699;
  wire seg_10_12_local_g2_3_42700;
  wire seg_10_12_local_g2_5_42702;
  wire seg_10_12_local_g2_6_42703;
  wire seg_10_12_local_g3_3_42708;
  wire seg_10_12_lutff_1_out_38810;
  wire seg_10_12_lutff_5_out_38814;
  wire seg_10_12_lutff_7_out_38816;
  wire seg_10_12_neigh_op_bot_0_38686;
  wire seg_10_12_neigh_op_bot_1_38687;
  wire seg_10_12_neigh_op_bot_4_38690;
  wire seg_10_12_neigh_op_rgt_6_42646;
  wire seg_10_12_sp4_h_r_11_42778;
  wire seg_10_12_sp4_h_r_12_38945;
  wire seg_10_12_sp4_h_r_16_38951;
  wire seg_10_12_sp4_h_r_35_35116;
  wire seg_10_12_sp4_h_r_4_42781;
  wire seg_10_12_sp4_h_r_6_42783;
  wire seg_10_12_sp4_h_r_8_42785;
  wire seg_10_12_sp4_r_v_b_27_42666;
  wire seg_10_12_sp4_r_v_b_35_42674;
  wire seg_10_12_sp4_v_b_13_38711;
  wire seg_10_12_sp4_v_b_17_38715;
  wire seg_10_12_sp4_v_b_1_38587;
  wire seg_10_12_sp4_v_b_20_38718;
  wire seg_10_12_sp4_v_b_22_38720;
  wire seg_10_12_sp4_v_b_23_38721;
  wire seg_10_12_sp4_v_b_25_38833;
  wire seg_10_12_sp4_v_b_34_38844;
  wire seg_10_12_sp4_v_b_45_38965;
  wire seg_10_13_glb_netwk_0_5;
  wire seg_10_13_local_g0_0_42804;
  wire seg_10_13_local_g0_1_42805;
  wire seg_10_13_local_g0_3_42807;
  wire seg_10_13_local_g0_4_42808;
  wire seg_10_13_local_g0_5_42809;
  wire seg_10_13_local_g0_6_42810;
  wire seg_10_13_local_g0_7_42811;
  wire seg_10_13_local_g1_0_42812;
  wire seg_10_13_local_g1_1_42813;
  wire seg_10_13_local_g1_3_42815;
  wire seg_10_13_local_g1_5_42817;
  wire seg_10_13_local_g2_2_42822;
  wire seg_10_13_local_g2_3_42823;
  wire seg_10_13_local_g3_0_42828;
  wire seg_10_13_local_g3_3_42831;
  wire seg_10_13_local_g3_4_42832;
  wire seg_10_13_local_g3_7_42835;
  wire seg_10_13_lutff_1_out_38933;
  wire seg_10_13_lutff_2_out_38934;
  wire seg_10_13_lutff_4_out_38936;
  wire seg_10_13_lutff_5_out_38937;
  wire seg_10_13_lutff_6_out_38938;
  wire seg_10_13_lutff_7_out_38939;
  wire seg_10_13_neigh_op_rgt_3_42766;
  wire seg_10_13_neigh_op_rgt_7_42770;
  wire seg_10_13_neigh_op_top_0_39055;
  wire seg_10_13_neigh_op_top_1_39056;
  wire seg_10_13_neigh_op_top_3_39058;
  wire seg_10_13_sp4_h_r_0_42898;
  wire seg_10_13_sp4_h_r_23_39069;
  wire seg_10_13_sp4_h_r_6_42906;
  wire seg_10_13_sp4_r_v_b_19_42671;
  wire seg_10_13_sp4_r_v_b_30_42794;
  wire seg_10_13_sp4_v_b_13_38834;
  wire seg_10_13_sp4_v_b_16_38837;
  wire seg_10_13_sp4_v_b_17_38838;
  wire seg_10_13_sp4_v_b_19_38840;
  wire seg_10_13_sp4_v_b_20_38841;
  wire seg_10_13_sp4_v_b_21_38842;
  wire seg_10_13_sp4_v_b_24_38957;
  wire seg_10_13_sp4_v_b_26_38959;
  wire seg_10_13_sp4_v_b_28_38961;
  wire seg_10_13_sp4_v_t_41_39207;
  wire seg_10_13_sp4_v_t_43_39209;
  wire seg_10_13_sp4_v_t_45_39211;
  wire seg_10_13_sp4_v_t_47_39213;
  wire seg_10_14_glb_netwk_0_5;
  wire seg_10_14_glb_netwk_1_6;
  wire seg_10_14_local_g0_0_42927;
  wire seg_10_14_local_g1_1_42936;
  wire seg_10_14_local_g1_3_42938;
  wire seg_10_14_local_g1_6_42941;
  wire seg_10_14_local_g1_7_42942;
  wire seg_10_14_local_g2_2_42945;
  wire seg_10_14_local_g2_4_42947;
  wire seg_10_14_local_g3_7_42958;
  wire seg_10_14_lutff_0_out_39055;
  wire seg_10_14_lutff_1_out_39056;
  wire seg_10_14_lutff_2_out_39057;
  wire seg_10_14_lutff_3_out_39058;
  wire seg_10_14_lutff_4_out_39059;
  wire seg_10_14_lutff_6_out_39061;
  wire seg_10_14_lutff_7_out_39062;
  wire seg_10_14_sp4_h_r_4_43027;
  wire seg_10_14_sp4_h_r_7_43030;
  wire seg_10_14_sp4_h_r_8_43031;
  wire seg_10_14_sp4_h_r_9_43032;
  wire seg_10_14_sp4_r_v_b_11_42674;
  wire seg_10_14_sp4_r_v_b_3_42666;
  wire seg_10_14_sp4_v_b_11_38843;
  wire seg_10_14_sp4_v_t_36_39325;
  wire seg_10_14_sp4_v_t_37_39326;
  wire seg_10_14_sp4_v_t_38_39327;
  wire seg_10_14_sp4_v_t_39_39328;
  wire seg_10_14_sp4_v_t_41_39330;
  wire seg_10_14_sp4_v_t_43_39332;
  wire seg_10_14_sp4_v_t_45_39334;
  wire seg_10_14_sp4_v_t_47_39336;
  wire seg_10_15_glb_netwk_0_5;
  wire seg_10_15_glb_netwk_1_6;
  wire seg_10_15_local_g0_2_43052;
  wire seg_10_15_local_g0_6_43056;
  wire seg_10_15_local_g3_0_43074;
  wire seg_10_15_lutff_2_out_39180;
  wire seg_10_15_sp4_h_r_4_43150;
  wire seg_10_15_sp4_h_r_6_43152;
  wire seg_10_15_sp4_v_b_0_38957;
  wire seg_10_15_sp4_v_b_32_39211;
  wire seg_10_15_sp4_v_b_8_38965;
  wire seg_10_15_sp4_v_t_36_39448;
  wire seg_10_15_sp4_v_t_43_39455;
  wire seg_10_16_sp4_v_b_1_39079;
  wire seg_10_16_sp4_v_t_42_39577;
  wire seg_10_16_sp4_v_t_44_39579;
  wire seg_10_17_glb_netwk_0_5;
  wire seg_10_17_local_g0_4_43300;
  wire seg_10_17_local_g0_6_43302;
  wire seg_10_17_local_g1_5_43309;
  wire seg_10_17_local_g1_7_43311;
  wire seg_10_17_local_g2_3_43315;
  wire seg_10_17_local_g3_1_43321;
  wire seg_10_17_local_g3_2_43322;
  wire seg_10_17_local_g3_5_43325;
  wire seg_10_17_lutff_2_out_39426;
  wire seg_10_17_lutff_3_out_39427;
  wire seg_10_17_lutff_4_out_39428;
  wire seg_10_17_lutff_5_out_39429;
  wire seg_10_17_lutff_6_out_39430;
  wire seg_10_17_lutff_7_out_39431;
  wire seg_10_17_neigh_op_bnr_5_43137;
  wire seg_10_17_neigh_op_rgt_1_43256;
  wire seg_10_17_sp4_h_l_39_28343;
  wire seg_10_17_sp4_h_r_14_39564;
  wire seg_10_17_sp4_h_r_20_39570;
  wire seg_10_17_sp4_h_r_26_35732;
  wire seg_10_17_sp4_h_r_28_35734;
  wire seg_10_17_sp4_h_r_6_43398;
  wire seg_10_17_sp4_h_r_8_43400;
  wire seg_10_17_sp4_r_v_b_11_43043;
  wire seg_10_17_sp4_r_v_b_13_43157;
  wire seg_10_17_sp4_r_v_b_15_43159;
  wire seg_10_17_sp4_r_v_b_25_43279;
  wire seg_10_17_sp4_r_v_b_27_43281;
  wire seg_10_17_sp4_r_v_b_29_43283;
  wire seg_10_17_sp4_r_v_b_31_43285;
  wire seg_10_17_sp4_r_v_b_37_43403;
  wire seg_10_17_sp4_r_v_b_39_43405;
  wire seg_10_17_sp4_r_v_b_41_43407;
  wire seg_10_17_sp4_r_v_b_5_43037;
  wire seg_10_17_sp4_r_v_b_9_43041;
  wire seg_10_17_sp4_v_b_10_39213;
  wire seg_10_17_sp4_v_b_12_39325;
  wire seg_10_17_sp4_v_b_14_39327;
  wire seg_10_17_sp4_v_b_30_39455;
  wire seg_10_17_sp4_v_b_42_39577;
  wire seg_10_17_sp4_v_b_44_39579;
  wire seg_10_17_sp4_v_b_4_39207;
  wire seg_10_17_sp4_v_b_6_39209;
  wire seg_10_17_sp4_v_b_8_39211;
  wire seg_10_18_glb_netwk_0_5;
  wire seg_10_18_local_g0_5_43424;
  wire seg_10_18_local_g1_3_43430;
  wire seg_10_18_local_g2_1_43436;
  wire seg_10_18_local_g2_2_43437;
  wire seg_10_18_local_g2_6_43441;
  wire seg_10_18_local_g3_0_43443;
  wire seg_10_18_local_g3_4_43447;
  wire seg_10_18_local_g3_7_43450;
  wire seg_10_18_lutff_0_out_39547;
  wire seg_10_18_lutff_1_out_39548;
  wire seg_10_18_lutff_2_out_39549;
  wire seg_10_18_lutff_3_out_39550;
  wire seg_10_18_lutff_4_out_39551;
  wire seg_10_18_lutff_5_out_39552;
  wire seg_10_18_lutff_6_out_39553;
  wire seg_10_18_lutff_7_out_39554;
  wire seg_10_18_sp4_h_r_14_39687;
  wire seg_10_18_sp4_h_r_16_39689;
  wire seg_10_18_sp4_h_r_18_39691;
  wire seg_10_18_sp4_h_r_22_39685;
  wire seg_10_18_sp4_h_r_24_35851;
  wire seg_10_18_sp4_h_r_26_35855;
  wire seg_10_18_sp4_h_r_32_35861;
  wire seg_10_18_sp4_h_r_34_35853;
  wire seg_10_18_sp4_h_r_4_43519;
  wire seg_10_18_sp4_h_r_8_43523;
  wire seg_10_18_sp4_r_v_b_11_43166;
  wire seg_10_18_sp4_r_v_b_13_43280;
  wire seg_10_18_sp4_r_v_b_15_43282;
  wire seg_10_18_sp4_r_v_b_19_43286;
  wire seg_10_18_sp4_r_v_b_1_43156;
  wire seg_10_18_sp4_r_v_b_23_43290;
  wire seg_10_18_sp4_r_v_b_31_43408;
  wire seg_10_18_sp4_r_v_b_37_43526;
  wire seg_10_18_sp4_r_v_b_39_43528;
  wire seg_10_18_sp4_r_v_b_3_43158;
  wire seg_10_18_sp4_r_v_b_43_43532;
  wire seg_10_18_sp4_r_v_b_45_43534;
  wire seg_10_18_sp4_r_v_b_5_43160;
  wire seg_10_18_sp4_r_v_b_9_43164;
  wire seg_10_18_sp4_v_b_0_39326;
  wire seg_10_18_sp4_v_b_10_39336;
  wire seg_10_18_sp4_v_b_11_39335;
  wire seg_10_18_sp4_v_b_12_39448;
  wire seg_10_18_sp4_v_b_2_39328;
  wire seg_10_18_sp4_v_b_4_39330;
  wire seg_10_18_sp4_v_b_6_39332;
  wire seg_10_18_sp4_v_b_7_39331;
  wire seg_10_18_sp4_v_b_8_39334;
  wire seg_10_19_glb_netwk_0_5;
  wire seg_10_19_local_g0_2_43544;
  wire seg_10_19_local_g0_6_43548;
  wire seg_10_19_local_g0_7_43549;
  wire seg_10_19_local_g1_0_43550;
  wire seg_10_19_local_g1_1_43551;
  wire seg_10_19_local_g1_4_43554;
  wire seg_10_19_local_g3_3_43569;
  wire seg_10_19_local_g3_5_43571;
  wire seg_10_19_lutff_0_out_39670;
  wire seg_10_19_lutff_1_out_39671;
  wire seg_10_19_lutff_2_out_39672;
  wire seg_10_19_lutff_3_out_39673;
  wire seg_10_19_lutff_4_out_39674;
  wire seg_10_19_lutff_5_out_39675;
  wire seg_10_19_lutff_6_out_39676;
  wire seg_10_19_lutff_7_out_39677;
  wire seg_10_19_sp4_h_r_0_43636;
  wire seg_10_19_sp4_h_r_10_43638;
  wire seg_10_19_sp4_h_r_12_39806;
  wire seg_10_19_sp4_h_r_14_39810;
  wire seg_10_19_sp4_h_r_16_39812;
  wire seg_10_19_sp4_h_r_20_39816;
  wire seg_10_19_sp4_h_r_24_35974;
  wire seg_10_19_sp4_h_r_28_35980;
  wire seg_10_19_sp4_h_r_2_43640;
  wire seg_10_19_sp4_h_r_34_35976;
  wire seg_10_19_sp4_h_r_4_43642;
  wire seg_10_19_sp4_h_r_6_43644;
  wire seg_10_19_sp4_h_r_8_43646;
  wire seg_10_19_sp4_r_v_b_21_43411;
  wire seg_10_19_sp4_r_v_b_23_43413;
  wire seg_10_20_glb_netwk_0_5;
  wire seg_10_20_local_g0_1_43666;
  wire seg_10_20_local_g0_3_43668;
  wire seg_10_20_local_g1_0_43673;
  wire seg_10_20_local_g3_2_43691;
  wire seg_10_20_lutff_0_out_39793;
  wire seg_10_20_lutff_1_out_39794;
  wire seg_10_20_lutff_2_out_39795;
  wire seg_10_20_lutff_3_out_39796;
  wire seg_10_20_sp12_h_r_12_21400;
  wire seg_10_20_sp4_h_r_0_43759;
  wire seg_10_20_sp4_h_r_22_39931;
  wire seg_10_20_sp4_h_r_2_43763;
  wire seg_10_20_sp4_h_r_4_43765;
  wire seg_10_20_sp4_h_r_6_43767;
  wire seg_10_20_sp4_v_b_1_39571;
  wire seg_10_21_sp4_v_b_2_39697;
  wire seg_10_22_sp4_v_b_10_39828;
  wire seg_10_24_sp4_v_b_9_40071;
  wire seg_10_25_sp4_v_b_10_40197;
  wire seg_10_26_glb_netwk_0_5;
  wire seg_10_26_local_g1_2_44413;
  wire seg_10_26_local_g3_3_44430;
  wire seg_10_26_local_g3_7_44434;
  wire seg_10_26_lutff_7_out_40538;
  wire seg_10_26_sp12_v_b_20_44250;
  wire seg_10_26_sp4_v_b_10_40320;
  wire seg_10_26_sp4_v_b_43_40685;
  wire seg_10_27_glb_netwk_0_5;
  wire seg_10_27_local_g0_3_44529;
  wire seg_10_27_local_g0_5_44531;
  wire seg_10_27_local_g0_6_44532;
  wire seg_10_27_local_g0_7_44533;
  wire seg_10_27_local_g1_3_44537;
  wire seg_10_27_local_g1_5_44539;
  wire seg_10_27_local_g1_7_44541;
  wire seg_10_27_local_g2_7_44549;
  wire seg_10_27_local_g3_3_44553;
  wire seg_10_27_local_g3_4_44554;
  wire seg_10_27_lutff_2_out_40656;
  wire seg_10_27_lutff_3_out_40657;
  wire seg_10_27_lutff_4_out_40658;
  wire seg_10_27_lutff_5_out_40659;
  wire seg_10_27_lutff_6_out_40660;
  wire seg_10_27_lutff_7_out_40661;
  wire seg_10_27_neigh_op_lft_5_36828;
  wire seg_10_27_neigh_op_lft_7_36830;
  wire seg_10_27_neigh_op_top_3_40780;
  wire seg_10_27_neigh_op_top_7_40784;
  wire seg_10_27_sp4_v_b_27_40680;
  wire seg_10_27_sp4_v_b_36_40801;
  wire seg_10_28_glb_netwk_0_5;
  wire seg_10_28_local_g0_4_44653;
  wire seg_10_28_local_g0_6_44655;
  wire seg_10_28_local_g0_7_44656;
  wire seg_10_28_local_g1_3_44660;
  wire seg_10_28_local_g1_6_44663;
  wire seg_10_28_local_g1_7_44664;
  wire seg_10_28_local_g2_5_44670;
  wire seg_10_28_local_g3_2_44675;
  wire seg_10_28_local_g3_3_44676;
  wire seg_10_28_local_g3_7_44680;
  wire seg_10_28_lutff_2_out_40779;
  wire seg_10_28_lutff_3_out_40780;
  wire seg_10_28_lutff_7_out_40784;
  wire seg_10_28_neigh_op_bnl_5_36828;
  wire seg_10_28_neigh_op_bnl_7_36830;
  wire seg_10_28_neigh_op_bot_4_40658;
  wire seg_10_28_neigh_op_bot_6_40660;
  wire seg_10_28_neigh_op_bot_7_40661;
  wire seg_10_28_neigh_op_tnl_3_37072;
  wire seg_10_28_neigh_op_top_6_40906;
  wire seg_10_28_sp4_v_b_26_40804;
  wire seg_10_29_glb_netwk_0_5;
  wire seg_10_29_local_g0_1_44773;
  wire seg_10_29_local_g0_2_44774;
  wire seg_10_29_local_g1_3_44783;
  wire seg_10_29_local_g1_4_44784;
  wire seg_10_29_local_g2_0_44788;
  wire seg_10_29_local_g2_5_44793;
  wire seg_10_29_local_g3_7_44803;
  wire seg_10_29_lutff_0_out_40900;
  wire seg_10_29_lutff_2_out_40902;
  wire seg_10_29_lutff_3_out_40903;
  wire seg_10_29_lutff_5_out_40905;
  wire seg_10_29_lutff_6_out_40906;
  wire seg_10_29_lutff_7_out_40907;
  wire seg_10_29_neigh_op_top_3_41026;
  wire seg_10_29_neigh_op_top_4_41027;
  wire seg_10_29_sp4_h_l_38_29568;
  wire seg_10_29_sp4_v_b_12_40801;
  wire seg_10_29_sp4_v_b_1_40678;
  wire seg_10_2_glb_netwk_0_5;
  wire seg_10_2_local_g0_2_41453;
  wire seg_10_2_local_g0_3_41454;
  wire seg_10_2_local_g0_4_41455;
  wire seg_10_2_local_g0_6_41457;
  wire seg_10_2_local_g0_7_41458;
  wire seg_10_2_local_g1_3_41462;
  wire seg_10_2_local_g1_4_41463;
  wire seg_10_2_local_g1_6_41465;
  wire seg_10_2_local_g2_4_41471;
  wire seg_10_2_local_g3_2_41477;
  wire seg_10_2_lutff_2_out_37545;
  wire seg_10_2_lutff_3_out_37546;
  wire seg_10_2_lutff_4_out_37547;
  wire seg_10_2_lutff_5_out_37548;
  wire seg_10_2_lutff_6_out_37549;
  wire seg_10_2_lutff_7_out_37550;
  wire seg_10_2_neigh_op_lft_4_33716;
  wire seg_10_2_neigh_op_top_2_37704;
  wire seg_10_2_neigh_op_top_3_37705;
  wire seg_10_2_neigh_op_top_4_37706;
  wire seg_10_2_neigh_op_top_6_37708;
  wire seg_10_2_sp4_v_b_19_37591;
  wire seg_10_30_glb_netwk_0_5;
  wire seg_10_30_local_g0_0_44895;
  wire seg_10_30_local_g0_2_44897;
  wire seg_10_30_local_g0_4_44899;
  wire seg_10_30_local_g0_5_44900;
  wire seg_10_30_local_g1_0_44903;
  wire seg_10_30_local_g1_2_44905;
  wire seg_10_30_local_g1_4_44907;
  wire seg_10_30_local_g1_5_44908;
  wire seg_10_30_local_g2_0_44911;
  wire seg_10_30_local_g2_2_44913;
  wire seg_10_30_local_g2_6_44917;
  wire seg_10_30_local_g3_3_44922;
  wire seg_10_30_local_g3_4_44923;
  wire seg_10_30_local_g3_6_44925;
  wire seg_10_30_local_g3_7_44926;
  wire seg_10_30_lutff_0_out_41023;
  wire seg_10_30_lutff_2_out_41025;
  wire seg_10_30_lutff_3_out_41026;
  wire seg_10_30_lutff_4_out_41027;
  wire seg_10_30_lutff_6_out_41029;
  wire seg_10_30_lutff_7_out_41030;
  wire seg_10_30_neigh_op_bot_0_40900;
  wire seg_10_30_neigh_op_bot_2_40902;
  wire seg_10_30_neigh_op_bot_5_40905;
  wire seg_10_30_neigh_op_lft_5_37197;
  wire seg_10_30_sp12_v_b_12_44250;
  wire seg_10_30_sp4_h_r_30_37331;
  wire seg_10_30_sp4_r_v_b_24_44879;
  wire seg_10_30_sp4_v_b_2_40804;
  wire seg_10_3_glb_netwk_0_5;
  wire seg_10_3_local_g0_2_41576;
  wire seg_10_3_local_g1_3_41585;
  wire seg_10_3_local_g1_5_41587;
  wire seg_10_3_local_g1_6_41588;
  wire seg_10_3_local_g2_4_41594;
  wire seg_10_3_local_g3_2_41600;
  wire seg_10_3_local_g3_3_41601;
  wire seg_10_3_local_g3_7_41605;
  wire seg_10_3_lutff_2_out_37704;
  wire seg_10_3_lutff_3_out_37705;
  wire seg_10_3_lutff_4_out_37706;
  wire seg_10_3_lutff_6_out_37708;
  wire seg_10_3_lutff_7_out_37709;
  wire seg_10_3_neigh_op_bnl_4_33716;
  wire seg_10_3_neigh_op_bot_3_37546;
  wire seg_10_3_neigh_op_bot_5_37548;
  wire seg_10_3_sp4_h_l_39_26915;
  wire seg_10_3_sp4_h_l_43_26919;
  wire seg_10_3_sp4_h_r_2_41672;
  wire seg_10_3_sp4_r_v_b_18_41435;
  wire seg_10_4_sp4_h_l_47_27015;
  wire seg_10_4_sp4_v_t_46_38105;
  wire seg_10_6_sp4_v_b_10_37860;
  wire seg_10_7_local_g0_5_42071;
  wire seg_10_7_local_g2_0_42082;
  wire seg_10_7_sp4_h_r_10_42162;
  wire seg_10_7_sp4_h_r_24_34498;
  wire seg_10_7_sp4_h_r_5_42167;
  wire seg_10_7_sp4_r_v_b_11_41813;
  wire seg_10_7_sp4_r_v_b_27_42051;
  wire seg_10_7_sp4_v_b_10_37983;
  wire seg_10_7_sp4_v_b_2_37975;
  wire seg_10_8_glb_netwk_0_5;
  wire seg_10_8_local_g0_3_42192;
  wire seg_10_8_local_g0_5_42194;
  wire seg_10_8_local_g0_6_42195;
  wire seg_10_8_local_g0_7_42196;
  wire seg_10_8_local_g1_0_42197;
  wire seg_10_8_local_g1_3_42200;
  wire seg_10_8_local_g1_6_42203;
  wire seg_10_8_local_g2_0_42205;
  wire seg_10_8_local_g2_4_42209;
  wire seg_10_8_local_g2_5_42210;
  wire seg_10_8_local_g2_6_42211;
  wire seg_10_8_local_g2_7_42212;
  wire seg_10_8_local_g3_3_42216;
  wire seg_10_8_local_g3_7_42220;
  wire seg_10_8_lutff_0_out_38317;
  wire seg_10_8_lutff_2_out_38319;
  wire seg_10_8_lutff_3_out_38320;
  wire seg_10_8_lutff_4_out_38321;
  wire seg_10_8_lutff_6_out_38323;
  wire seg_10_8_lutff_7_out_38324;
  wire seg_10_8_neigh_op_bnr_0_42025;
  wire seg_10_8_neigh_op_lft_5_34491;
  wire seg_10_8_neigh_op_lft_6_34492;
  wire seg_10_8_neigh_op_lft_7_34493;
  wire seg_10_8_neigh_op_rgt_5_42153;
  wire seg_10_8_neigh_op_rgt_6_42154;
  wire seg_10_8_neigh_op_rgt_7_42155;
  wire seg_10_8_sp4_r_v_b_30_42179;
  wire seg_10_8_sp4_r_v_b_32_42181;
  wire seg_10_8_sp4_r_v_b_35_42182;
  wire seg_10_8_sp4_r_v_b_36_42295;
  wire seg_10_8_sp4_v_b_10_38106;
  wire seg_10_8_sp4_v_b_43_38471;
  wire seg_10_8_sp4_v_t_38_38589;
  wire seg_10_9_sp4_h_r_11_42409;
  wire seg_10_9_sp4_h_r_5_42413;
  wire seg_10_9_sp4_v_b_10_38229;
  wire seg_10_9_sp4_v_b_8_38227;
  wire seg_11_10_glb_netwk_0_5;
  wire seg_11_10_local_g0_2_46268;
  wire seg_11_10_local_g0_3_46269;
  wire seg_11_10_local_g0_5_46271;
  wire seg_11_10_local_g0_7_46273;
  wire seg_11_10_local_g1_2_46276;
  wire seg_11_10_local_g1_3_46277;
  wire seg_11_10_local_g1_5_46279;
  wire seg_11_10_local_g2_4_46286;
  wire seg_11_10_local_g3_2_46292;
  wire seg_11_10_local_g3_4_46294;
  wire seg_11_10_local_g3_7_46297;
  wire seg_11_10_lutff_4_out_42398;
  wire seg_11_10_lutff_5_out_42399;
  wire seg_11_10_lutff_6_out_42400;
  wire seg_11_10_lutff_7_out_42401;
  wire seg_11_10_neigh_op_bot_7_42278;
  wire seg_11_10_sp4_h_l_36_31037;
  wire seg_11_10_sp4_h_r_11_46363;
  wire seg_11_10_sp4_h_r_12_42530;
  wire seg_11_10_sp4_h_r_13_42529;
  wire seg_11_10_sp4_h_r_14_42534;
  wire seg_11_10_sp4_h_r_24_38698;
  wire seg_11_10_sp4_h_r_26_38702;
  wire seg_11_10_sp4_h_r_36_34868;
  wire seg_11_10_sp4_h_r_3_46365;
  wire seg_11_10_sp4_h_r_6_46368;
  wire seg_11_10_sp4_h_r_8_46370;
  wire seg_11_10_sp4_r_v_b_13_46127;
  wire seg_11_10_sp4_r_v_b_25_46249;
  wire seg_11_10_sp4_r_v_b_26_46252;
  wire seg_11_10_sp4_r_v_b_29_46253;
  wire seg_11_10_sp4_r_v_b_31_46255;
  wire seg_11_10_sp4_r_v_b_33_46257;
  wire seg_11_10_sp4_r_v_b_39_46375;
  wire seg_11_10_sp4_r_v_b_41_46377;
  wire seg_11_10_sp4_r_v_b_47_46383;
  wire seg_11_10_sp4_r_v_b_9_46011;
  wire seg_11_10_sp4_v_b_11_42182;
  wire seg_11_10_sp4_v_b_12_42295;
  wire seg_11_10_sp4_v_b_24_42419;
  wire seg_11_10_sp4_v_b_40_42545;
  wire seg_11_10_sp4_v_b_44_42549;
  wire seg_11_11_glb_netwk_0_5;
  wire seg_11_11_glb_netwk_1_6;
  wire seg_11_11_local_g2_2_46407;
  wire seg_11_11_local_g3_6_46419;
  wire seg_11_11_lutff_2_out_42519;
  wire seg_11_11_lutff_7_out_42524;
  wire seg_11_11_sp4_r_v_b_22_46259;
  wire seg_11_11_sp4_v_b_26_42544;
  wire seg_11_11_sp4_v_t_46_42797;
  wire seg_11_12_glb_netwk_0_5;
  wire seg_11_12_glb_netwk_1_6;
  wire seg_11_12_local_g0_1_46513;
  wire seg_11_12_local_g0_2_46514;
  wire seg_11_12_local_g0_5_46517;
  wire seg_11_12_local_g0_7_46519;
  wire seg_11_12_local_g1_5_46525;
  wire seg_11_12_local_g2_1_46529;
  wire seg_11_12_local_g2_4_46532;
  wire seg_11_12_local_g2_5_46533;
  wire seg_11_12_local_g2_6_46534;
  wire seg_11_12_local_g2_7_46535;
  wire seg_11_12_local_g3_1_46537;
  wire seg_11_12_lutff_2_out_42642;
  wire seg_11_12_lutff_6_out_42646;
  wire seg_11_12_lutff_7_out_42647;
  wire seg_11_12_neigh_op_lft_1_38810;
  wire seg_11_12_neigh_op_lft_5_38814;
  wire seg_11_12_neigh_op_lft_7_38816;
  wire seg_11_12_neigh_op_rgt_1_46472;
  wire seg_11_12_neigh_op_rgt_5_46476;
  wire seg_11_12_neigh_op_rgt_7_46478;
  wire seg_11_12_sp4_h_r_14_42780;
  wire seg_11_12_sp4_h_r_20_42786;
  wire seg_11_12_sp4_h_r_2_46610;
  wire seg_11_12_sp4_h_r_6_46614;
  wire seg_11_12_sp4_h_r_8_46616;
  wire seg_11_12_sp4_r_v_b_14_46374;
  wire seg_11_12_sp4_r_v_b_17_46377;
  wire seg_11_12_sp4_v_b_0_42419;
  wire seg_11_12_sp4_v_b_21_42550;
  wire seg_11_12_sp4_v_b_28_42669;
  wire seg_11_12_sp4_v_t_41_42915;
  wire seg_11_12_sp4_v_t_45_42919;
  wire seg_11_12_sp4_v_t_47_42921;
  wire seg_11_13_local_g0_4_46639;
  wire seg_11_13_local_g0_5_46640;
  wire seg_11_13_local_g0_6_46641;
  wire seg_11_13_local_g0_7_46642;
  wire seg_11_13_local_g1_1_46644;
  wire seg_11_13_local_g1_2_46645;
  wire seg_11_13_local_g1_3_46646;
  wire seg_11_13_local_g1_4_46647;
  wire seg_11_13_local_g1_5_46648;
  wire seg_11_13_local_g1_7_46650;
  wire seg_11_13_local_g2_1_46652;
  wire seg_11_13_local_g2_2_46653;
  wire seg_11_13_local_g2_5_46656;
  wire seg_11_13_local_g2_7_46658;
  wire seg_11_13_local_g3_4_46663;
  wire seg_11_13_local_g3_6_46665;
  wire seg_11_13_lutff_3_out_42766;
  wire seg_11_13_lutff_7_out_42770;
  wire seg_11_13_neigh_op_bot_7_42647;
  wire seg_11_13_neigh_op_lft_1_38933;
  wire seg_11_13_neigh_op_lft_2_38934;
  wire seg_11_13_neigh_op_lft_4_38936;
  wire seg_11_13_neigh_op_lft_5_38937;
  wire seg_11_13_neigh_op_lft_6_38938;
  wire seg_11_13_neigh_op_lft_7_38939;
  wire seg_11_13_neigh_op_rgt_1_46595;
  wire seg_11_13_neigh_op_rgt_2_46596;
  wire seg_11_13_neigh_op_rgt_4_46598;
  wire seg_11_13_neigh_op_rgt_5_46599;
  wire seg_11_13_neigh_op_rgt_6_46600;
  wire seg_11_13_neigh_op_rgt_7_46601;
  wire seg_11_13_sp12_h_r_2_42895;
  wire seg_11_13_sp4_h_r_12_42899;
  wire seg_11_13_sp4_h_r_20_42909;
  wire seg_11_13_sp4_h_r_24_39067;
  wire seg_11_13_sp4_h_r_2_46733;
  wire seg_11_13_sp4_h_r_32_39077;
  wire seg_11_13_sp4_h_r_4_46735;
  wire seg_11_13_sp4_r_v_b_3_46374;
  wire seg_11_13_sp4_v_b_5_42545;
  wire seg_11_13_sp4_v_b_9_42549;
  wire seg_11_13_sp4_v_t_37_43034;
  wire seg_11_13_sp4_v_t_39_43036;
  wire seg_11_13_sp4_v_t_40_43037;
  wire seg_11_13_sp4_v_t_44_43041;
  wire seg_11_13_sp4_v_t_45_43042;
  wire seg_11_13_sp4_v_t_46_43043;
  wire seg_11_14_glb_netwk_0_5;
  wire seg_11_14_local_g0_0_46758;
  wire seg_11_14_local_g0_2_46760;
  wire seg_11_14_local_g0_4_46762;
  wire seg_11_14_local_g0_6_46764;
  wire seg_11_14_local_g0_7_46765;
  wire seg_11_14_local_g1_2_46768;
  wire seg_11_14_local_g1_3_46769;
  wire seg_11_14_local_g1_7_46773;
  wire seg_11_14_local_g2_0_46774;
  wire seg_11_14_local_g2_2_46776;
  wire seg_11_14_local_g2_6_46780;
  wire seg_11_14_local_g3_2_46784;
  wire seg_11_14_lutff_0_out_42886;
  wire seg_11_14_lutff_2_out_42888;
  wire seg_11_14_lutff_3_out_42889;
  wire seg_11_14_lutff_4_out_42890;
  wire seg_11_14_lutff_6_out_42892;
  wire seg_11_14_neigh_op_lft_4_39059;
  wire seg_11_14_neigh_op_lft_6_39061;
  wire seg_11_14_neigh_op_lft_7_39062;
  wire seg_11_14_sp4_h_r_10_46854;
  wire seg_11_14_sp4_h_r_14_43026;
  wire seg_11_14_sp4_h_r_2_46856;
  wire seg_11_14_sp4_h_r_34_39192;
  wire seg_11_14_sp4_h_r_7_46861;
  wire seg_11_14_sp4_h_r_8_46862;
  wire seg_11_14_sp4_r_v_b_27_46743;
  wire seg_11_14_sp4_r_v_b_3_46497;
  wire seg_11_14_sp4_r_v_b_42_46870;
  wire seg_11_14_sp4_v_b_0_42665;
  wire seg_11_14_sp4_v_b_2_42667;
  wire seg_11_14_sp4_v_t_36_43156;
  wire seg_11_14_sp4_v_t_37_43157;
  wire seg_11_14_sp4_v_t_38_43158;
  wire seg_11_14_sp4_v_t_39_43159;
  wire seg_11_14_sp4_v_t_40_43160;
  wire seg_11_14_sp4_v_t_42_43162;
  wire seg_11_14_sp4_v_t_44_43164;
  wire seg_11_14_sp4_v_t_46_43166;
  wire seg_11_15_glb_netwk_0_5;
  wire seg_11_15_local_g0_3_46884;
  wire seg_11_15_local_g1_3_46892;
  wire seg_11_15_local_g1_5_46894;
  wire seg_11_15_local_g2_1_46898;
  wire seg_11_15_local_g3_0_46905;
  wire seg_11_15_lutff_2_out_43011;
  wire seg_11_15_lutff_4_out_43013;
  wire seg_11_15_lutff_6_out_43015;
  wire seg_11_15_neigh_op_rgt_0_46840;
  wire seg_11_15_sp4_h_r_3_46980;
  wire seg_11_15_sp4_h_r_5_46982;
  wire seg_11_15_sp4_r_v_b_27_46866;
  wire seg_11_15_sp4_v_b_33_43041;
  wire seg_11_15_sp4_v_b_6_42794;
  wire seg_11_15_sp4_v_t_36_43279;
  wire seg_11_15_sp4_v_t_37_43280;
  wire seg_11_15_sp4_v_t_38_43281;
  wire seg_11_15_sp4_v_t_40_43283;
  wire seg_11_15_sp4_v_t_42_43285;
  wire seg_11_15_sp4_v_t_43_43286;
  wire seg_11_15_sp4_v_t_47_43290;
  wire seg_11_16_glb_netwk_0_5;
  wire seg_11_16_local_g0_2_47006;
  wire seg_11_16_local_g0_5_47009;
  wire seg_11_16_lutff_5_out_43137;
  wire seg_11_16_sp4_h_r_10_47100;
  wire seg_11_16_sp4_r_v_b_11_46751;
  wire seg_11_16_sp4_r_v_b_43_47117;
  wire seg_11_16_sp4_v_b_18_43039;
  wire seg_11_16_sp4_v_t_37_43403;
  wire seg_11_16_sp4_v_t_39_43405;
  wire seg_11_16_sp4_v_t_41_43407;
  wire seg_11_17_glb_netwk_0_5;
  wire seg_11_17_local_g0_1_47128;
  wire seg_11_17_local_g2_5_47148;
  wire seg_11_17_lutff_1_out_43256;
  wire seg_11_17_sp4_h_r_18_43399;
  wire seg_11_17_sp4_h_r_2_47225;
  wire seg_11_17_sp4_r_v_b_13_46988;
  wire seg_11_17_sp4_r_v_b_35_47120;
  wire seg_11_17_sp4_v_b_18_43162;
  wire seg_11_17_sp4_v_t_37_43526;
  wire seg_11_17_sp4_v_t_39_43528;
  wire seg_11_17_sp4_v_t_43_43532;
  wire seg_11_17_sp4_v_t_45_43534;
  wire seg_11_18_glb_netwk_0_5;
  wire seg_11_18_local_g0_2_47252;
  wire seg_11_18_local_g1_0_47258;
  wire seg_11_18_local_g2_2_47268;
  wire seg_11_18_local_g2_3_47269;
  wire seg_11_18_local_g2_5_47271;
  wire seg_11_18_local_g2_6_47272;
  wire seg_11_18_local_g3_0_47274;
  wire seg_11_18_local_g3_1_47275;
  wire seg_11_18_local_g3_2_47276;
  wire seg_11_18_local_g3_5_47279;
  wire seg_11_18_lutff_3_out_43381;
  wire seg_11_18_lutff_4_out_43382;
  wire seg_11_18_lutff_5_out_43383;
  wire seg_11_18_neigh_op_tnl_0_39670;
  wire seg_11_18_neigh_op_tnl_5_39675;
  wire seg_11_18_neigh_op_tnl_6_39676;
  wire seg_11_18_sp4_h_r_16_43520;
  wire seg_11_18_sp4_h_r_26_39686;
  wire seg_11_18_sp4_h_r_2_47348;
  wire seg_11_18_sp4_h_r_34_39684;
  wire seg_11_18_sp4_h_r_4_47350;
  wire seg_11_18_sp4_r_v_b_41_47361;
  wire seg_11_18_sp4_v_b_10_43167;
  wire seg_11_19_glb_netwk_0_5;
  wire seg_11_19_local_g0_1_47374;
  wire seg_11_19_local_g0_4_47377;
  wire seg_11_19_local_g1_1_47382;
  wire seg_11_19_local_g1_4_47385;
  wire seg_11_19_local_g2_2_47391;
  wire seg_11_19_local_g3_0_47397;
  wire seg_11_19_local_g3_6_47403;
  wire seg_11_19_lutff_2_out_43503;
  wire seg_11_19_lutff_6_out_43507;
  wire seg_11_19_neigh_op_lft_1_39671;
  wire seg_11_19_neigh_op_lft_4_39674;
  wire seg_11_19_neigh_op_top_1_43625;
  wire seg_11_19_sp4_h_r_6_47475;
  wire seg_11_19_sp4_r_v_b_16_47237;
  wire seg_11_19_sp4_r_v_b_28_47361;
  wire seg_11_19_sp4_v_b_2_43282;
  wire seg_11_19_sp4_v_b_34_43536;
  wire seg_11_20_glb_netwk_0_5;
  wire seg_11_20_glb_netwk_1_6;
  wire seg_11_20_local_g0_2_47498;
  wire seg_11_20_local_g1_1_47505;
  wire seg_11_20_local_g2_4_47516;
  wire seg_11_20_lutff_1_out_43625;
  wire seg_11_20_neigh_op_bnl_4_39674;
  wire seg_11_20_neigh_op_lft_1_39794;
  wire seg_11_20_neigh_op_lft_2_39795;
  wire seg_11_20_sp4_h_r_12_43760;
  wire seg_11_20_sp4_h_r_4_47596;
  wire seg_11_20_sp4_v_b_10_43413;
  wire seg_11_20_sp4_v_b_7_43408;
  wire seg_11_20_sp4_v_b_8_43411;
  wire seg_11_21_sp4_h_r_5_47720;
  wire seg_11_22_sp4_v_t_44_44148;
  wire seg_11_23_glb_netwk_0_5;
  wire seg_11_23_local_g2_2_47883;
  wire seg_11_23_local_g3_3_47892;
  wire seg_11_23_sp4_r_v_b_13_47726;
  wire seg_11_23_sp4_r_v_b_19_47732;
  wire seg_11_23_sp4_v_b_34_44028;
  wire seg_11_23_sp4_v_b_44_44148;
  wire seg_11_25_sp4_v_t_47_44520;
  wire seg_11_29_local_g0_3_48606;
  wire seg_11_29_local_g1_5_48616;
  wire seg_11_29_neigh_op_lft_3_40903;
  wire seg_11_29_neigh_op_lft_5_40905;
  wire seg_11_29_sp4_v_b_10_44520;
  wire seg_11_30_local_g1_3_48737;
  wire seg_11_30_local_g1_4_48738;
  wire seg_11_30_local_g2_0_48742;
  wire seg_11_30_local_g2_5_48747;
  wire seg_11_30_neigh_op_bnl_0_40900;
  wire seg_11_30_neigh_op_bnl_5_40905;
  wire seg_11_30_neigh_op_lft_3_41026;
  wire seg_11_30_neigh_op_lft_4_41027;
  wire seg_11_30_sp4_h_r_6_48824;
  wire seg_11_31_span4_horz_l_14_33556;
  wire seg_11_4_sp4_h_l_42_30307;
  wire seg_11_7_glb_netwk_0_5;
  wire seg_11_7_local_g1_2_45907;
  wire seg_11_7_local_g1_3_45908;
  wire seg_11_7_local_g1_6_45911;
  wire seg_11_7_local_g1_7_45912;
  wire seg_11_7_local_g3_0_45921;
  wire seg_11_7_local_g3_2_45923;
  wire seg_11_7_local_g3_3_45924;
  wire seg_11_7_lutff_0_out_42025;
  wire seg_11_7_lutff_2_out_42027;
  wire seg_11_7_lutff_7_out_42032;
  wire seg_11_7_sp4_h_r_6_45999;
  wire seg_11_7_sp4_r_v_b_17_45762;
  wire seg_11_7_sp4_r_v_b_18_45763;
  wire seg_11_7_sp4_v_b_11_41813;
  wire seg_11_7_sp4_v_b_43_42179;
  wire seg_11_7_sp4_v_t_36_42295;
  wire seg_11_8_local_g0_0_46020;
  wire seg_11_8_local_g0_1_46021;
  wire seg_11_8_local_g0_2_46022;
  wire seg_11_8_local_g0_3_46023;
  wire seg_11_8_local_g0_4_46024;
  wire seg_11_8_local_g1_0_46028;
  wire seg_11_8_local_g1_2_46030;
  wire seg_11_8_local_g1_6_46034;
  wire seg_11_8_local_g1_7_46035;
  wire seg_11_8_local_g2_1_46037;
  wire seg_11_8_lutff_2_out_42150;
  wire seg_11_8_lutff_3_out_42151;
  wire seg_11_8_lutff_4_out_42152;
  wire seg_11_8_lutff_5_out_42153;
  wire seg_11_8_lutff_6_out_42154;
  wire seg_11_8_lutff_7_out_42155;
  wire seg_11_8_neigh_op_bot_0_42025;
  wire seg_11_8_neigh_op_lft_2_38319;
  wire seg_11_8_neigh_op_lft_4_38321;
  wire seg_11_8_neigh_op_lft_6_38323;
  wire seg_11_8_neigh_op_rgt_1_45980;
  wire seg_11_8_neigh_op_top_0_42271;
  wire seg_11_8_neigh_op_top_1_42272;
  wire seg_11_8_neigh_op_top_3_42274;
  wire seg_11_8_sp4_h_l_37_30790;
  wire seg_11_8_sp4_r_v_b_2_45760;
  wire seg_11_8_sp4_r_v_b_7_45763;
  wire seg_11_8_sp4_v_b_0_41927;
  wire seg_11_9_glb_netwk_0_5;
  wire seg_11_9_local_g0_2_46145;
  wire seg_11_9_local_g0_3_46146;
  wire seg_11_9_local_g0_4_46147;
  wire seg_11_9_local_g0_5_46148;
  wire seg_11_9_local_g0_6_46149;
  wire seg_11_9_local_g0_7_46150;
  wire seg_11_9_local_g1_3_46154;
  wire seg_11_9_local_g1_4_46155;
  wire seg_11_9_local_g1_5_46156;
  wire seg_11_9_local_g1_6_46157;
  wire seg_11_9_local_g1_7_46158;
  wire seg_11_9_local_g2_6_46165;
  wire seg_11_9_local_g3_0_46167;
  wire seg_11_9_lutff_0_out_42271;
  wire seg_11_9_lutff_1_out_42272;
  wire seg_11_9_lutff_3_out_42274;
  wire seg_11_9_lutff_4_out_42275;
  wire seg_11_9_lutff_5_out_42276;
  wire seg_11_9_lutff_6_out_42277;
  wire seg_11_9_lutff_7_out_42278;
  wire seg_11_9_neigh_op_bnr_5_45984;
  wire seg_11_9_neigh_op_bot_2_42150;
  wire seg_11_9_neigh_op_bot_3_42151;
  wire seg_11_9_neigh_op_bot_4_42152;
  wire seg_11_9_neigh_op_top_6_42400;
  wire seg_11_9_sp4_h_r_15_42410;
  wire seg_11_9_sp4_h_r_16_42413;
  wire seg_11_9_sp4_h_r_22_42409;
  wire seg_11_9_sp4_h_r_23_42408;
  wire seg_11_9_sp4_h_r_34_38577;
  wire seg_11_9_sp4_v_b_14_42174;
  wire seg_11_9_sp4_v_b_3_42051;
  wire seg_11_9_sp4_v_b_40_42422;
  wire seg_12_0_local_g0_3_48895;
  wire seg_12_0_local_g0_3_48895_i1;
  wire seg_12_0_local_g0_3_48895_i2;
  wire seg_12_0_local_g0_3_48895_i3;
  wire seg_12_0_span4_vert_19_45240;
  wire seg_12_0_span4_vert_25_45247;
  wire seg_12_10_sp12_v_b_23_50067;
  wire seg_12_10_sp4_v_b_4_46008;
  wire seg_12_10_sp4_v_b_9_46011;
  wire seg_12_11_glb_netwk_0_5;
  wire seg_12_11_local_g0_0_50220;
  wire seg_12_11_local_g0_3_50223;
  wire seg_12_11_local_g0_6_50226;
  wire seg_12_11_local_g0_7_50227;
  wire seg_12_11_local_g1_1_50229;
  wire seg_12_11_local_g1_2_50230;
  wire seg_12_11_local_g1_6_50234;
  wire seg_12_11_local_g2_3_50239;
  wire seg_12_11_local_g2_4_50240;
  wire seg_12_11_local_g3_3_50247;
  wire seg_12_11_lutff_0_out_46348;
  wire seg_12_11_lutff_2_out_46350;
  wire seg_12_11_lutff_5_out_46353;
  wire seg_12_11_lutff_6_out_46354;
  wire seg_12_11_neigh_op_bnl_4_42398;
  wire seg_12_11_neigh_op_lft_2_42519;
  wire seg_12_11_neigh_op_lft_7_42524;
  wire seg_12_11_sp12_v_t_23_50313;
  wire seg_12_11_sp4_h_r_17_46489;
  wire seg_12_11_sp4_h_r_2_50318;
  wire seg_12_11_sp4_r_v_b_23_50091;
  wire seg_12_11_sp4_r_v_b_32_50212;
  wire seg_12_11_sp4_v_b_22_46259;
  wire seg_12_11_sp4_v_b_27_46374;
  wire seg_12_11_sp4_v_b_35_46382;
  wire seg_12_11_sp4_v_t_38_46620;
  wire seg_12_11_sp4_v_t_42_46624;
  wire seg_12_12_glb_netwk_0_5;
  wire seg_12_12_local_g0_0_50343;
  wire seg_12_12_local_g0_1_50344;
  wire seg_12_12_local_g0_2_50345;
  wire seg_12_12_local_g0_3_50346;
  wire seg_12_12_local_g0_4_50347;
  wire seg_12_12_local_g0_5_50348;
  wire seg_12_12_local_g0_6_50349;
  wire seg_12_12_local_g1_0_50351;
  wire seg_12_12_local_g1_2_50353;
  wire seg_12_12_local_g1_3_50354;
  wire seg_12_12_local_g1_4_50355;
  wire seg_12_12_local_g1_5_50356;
  wire seg_12_12_local_g2_0_50359;
  wire seg_12_12_local_g2_1_50360;
  wire seg_12_12_local_g2_2_50361;
  wire seg_12_12_local_g3_3_50370;
  wire seg_12_12_local_g3_4_50371;
  wire seg_12_12_lutff_1_out_46472;
  wire seg_12_12_lutff_3_out_46474;
  wire seg_12_12_lutff_4_out_46475;
  wire seg_12_12_lutff_5_out_46476;
  wire seg_12_12_lutff_6_out_46477;
  wire seg_12_12_lutff_7_out_46478;
  wire seg_12_12_neigh_op_bnr_1_50180;
  wire seg_12_12_neigh_op_bot_2_46350;
  wire seg_12_12_neigh_op_bot_5_46353;
  wire seg_12_12_neigh_op_rgt_4_50306;
  wire seg_12_12_sp4_h_r_11_50440;
  wire seg_12_12_sp4_h_r_12_46607;
  wire seg_12_12_sp4_h_r_14_46611;
  wire seg_12_12_sp4_h_r_16_46613;
  wire seg_12_12_sp4_h_r_18_46615;
  wire seg_12_12_sp4_h_r_20_46617;
  wire seg_12_12_sp4_h_r_2_50441;
  wire seg_12_12_sp4_h_r_4_50443;
  wire seg_12_12_sp4_r_v_b_33_50334;
  wire seg_12_12_sp4_v_b_10_46260;
  wire seg_12_12_sp4_v_b_13_46373;
  wire seg_12_12_sp4_v_b_16_46376;
  wire seg_12_12_sp4_v_b_19_46379;
  wire seg_12_12_sp4_v_b_1_46249;
  wire seg_12_12_sp4_v_b_32_46504;
  wire seg_12_12_sp4_v_b_42_46624;
  wire seg_12_12_sp4_v_b_43_46625;
  wire seg_12_12_sp4_v_b_5_46253;
  wire seg_12_12_sp4_v_b_7_46255;
  wire seg_12_12_sp4_v_t_46_46751;
  wire seg_12_13_glb_netwk_0_5;
  wire seg_12_13_local_g0_0_50466;
  wire seg_12_13_local_g0_1_50467;
  wire seg_12_13_local_g0_2_50468;
  wire seg_12_13_local_g0_3_50469;
  wire seg_12_13_local_g0_5_50471;
  wire seg_12_13_local_g1_0_50474;
  wire seg_12_13_local_g1_1_50475;
  wire seg_12_13_local_g1_3_50477;
  wire seg_12_13_local_g1_4_50478;
  wire seg_12_13_local_g1_5_50479;
  wire seg_12_13_local_g1_7_50481;
  wire seg_12_13_local_g2_1_50483;
  wire seg_12_13_local_g2_2_50484;
  wire seg_12_13_local_g2_3_50485;
  wire seg_12_13_local_g3_2_50492;
  wire seg_12_13_local_g3_3_50493;
  wire seg_12_13_local_g3_5_50495;
  wire seg_12_13_lutff_0_out_46594;
  wire seg_12_13_lutff_1_out_46595;
  wire seg_12_13_lutff_2_out_46596;
  wire seg_12_13_lutff_3_out_46597;
  wire seg_12_13_lutff_4_out_46598;
  wire seg_12_13_lutff_5_out_46599;
  wire seg_12_13_lutff_6_out_46600;
  wire seg_12_13_lutff_7_out_46601;
  wire seg_12_13_neigh_op_tnl_2_42888;
  wire seg_12_13_neigh_op_tnl_3_42889;
  wire seg_12_13_neigh_op_tnr_2_50550;
  wire seg_12_13_neigh_op_top_1_46718;
  wire seg_12_13_neigh_op_top_3_46720;
  wire seg_12_13_neigh_op_top_5_46722;
  wire seg_12_13_sp4_h_r_16_46736;
  wire seg_12_13_sp4_h_r_18_46738;
  wire seg_12_13_sp4_h_r_1_50561;
  wire seg_12_13_sp4_h_r_21_46739;
  wire seg_12_13_sp4_h_r_43_39075;
  wire seg_12_13_sp4_h_r_8_50570;
  wire seg_12_13_sp4_r_v_b_21_50335;
  wire seg_12_13_sp4_r_v_b_27_50451;
  wire seg_12_13_sp4_r_v_b_9_50211;
  wire seg_12_13_sp4_v_b_10_46383;
  wire seg_12_13_sp4_v_b_12_46495;
  wire seg_12_13_sp4_v_b_15_46498;
  wire seg_12_13_sp4_v_b_17_46500;
  wire seg_12_13_sp4_v_b_2_46375;
  wire seg_12_13_sp4_v_b_4_46377;
  wire seg_12_13_sp4_v_t_38_46866;
  wire seg_12_13_sp4_v_t_39_46867;
  wire seg_12_13_sp4_v_t_41_46869;
  wire seg_12_13_sp4_v_t_42_46870;
  wire seg_12_13_sp4_v_t_45_46873;
  wire seg_12_14_glb_netwk_0_5;
  wire seg_12_14_local_g0_4_50593;
  wire seg_12_14_local_g1_0_50597;
  wire seg_12_14_local_g1_1_50598;
  wire seg_12_14_local_g1_2_50599;
  wire seg_12_14_local_g1_3_50600;
  wire seg_12_14_local_g1_4_50601;
  wire seg_12_14_local_g1_5_50602;
  wire seg_12_14_local_g1_6_50603;
  wire seg_12_14_local_g2_4_50609;
  wire seg_12_14_local_g3_0_50613;
  wire seg_12_14_local_g3_2_50615;
  wire seg_12_14_local_g3_3_50616;
  wire seg_12_14_local_g3_4_50617;
  wire seg_12_14_local_g3_7_50620;
  wire seg_12_14_lutff_0_out_46717;
  wire seg_12_14_lutff_1_out_46718;
  wire seg_12_14_lutff_3_out_46720;
  wire seg_12_14_lutff_4_out_46721;
  wire seg_12_14_lutff_5_out_46722;
  wire seg_12_14_neigh_op_lft_4_42890;
  wire seg_12_14_neigh_op_rgt_7_50555;
  wire seg_12_14_neigh_op_tnl_4_43013;
  wire seg_12_14_sp4_h_r_10_50685;
  wire seg_12_14_sp4_h_r_14_46857;
  wire seg_12_14_sp4_h_r_19_46860;
  wire seg_12_14_sp4_h_r_28_43027;
  wire seg_12_14_sp4_h_r_4_50689;
  wire seg_12_14_sp4_r_v_b_2_50329;
  wire seg_12_14_sp4_r_v_b_30_50579;
  wire seg_12_14_sp4_r_v_b_40_50699;
  wire seg_12_14_sp4_r_v_b_5_50330;
  wire seg_12_14_sp4_v_b_0_46496;
  wire seg_12_14_sp4_v_b_42_46870;
  wire seg_12_14_sp4_v_b_43_46871;
  wire seg_12_14_sp4_v_b_8_46504;
  wire seg_12_14_sp4_v_b_9_46503;
  wire seg_12_14_sp4_v_t_36_46987;
  wire seg_12_14_sp4_v_t_43_46994;
  wire seg_12_14_sp4_v_t_45_46996;
  wire seg_12_14_sp4_v_t_47_46998;
  wire seg_12_15_glb_netwk_0_5;
  wire seg_12_15_glb_netwk_1_6;
  wire seg_12_15_local_g0_0_50712;
  wire seg_12_15_local_g0_1_50713;
  wire seg_12_15_local_g0_4_50716;
  wire seg_12_15_local_g0_6_50718;
  wire seg_12_15_local_g1_2_50722;
  wire seg_12_15_local_g1_4_50724;
  wire seg_12_15_local_g1_6_50726;
  wire seg_12_15_local_g2_0_50728;
  wire seg_12_15_local_g2_7_50735;
  wire seg_12_15_local_g3_4_50740;
  wire seg_12_15_local_g3_7_50743;
  wire seg_12_15_lutff_0_out_46840;
  wire seg_12_15_lutff_4_out_46844;
  wire seg_12_15_lutff_5_out_46845;
  wire seg_12_15_lutff_7_out_46847;
  wire seg_12_15_neigh_op_lft_2_43011;
  wire seg_12_15_neigh_op_lft_4_43013;
  wire seg_12_15_neigh_op_lft_6_43015;
  wire seg_12_15_sp4_h_r_14_46980;
  wire seg_12_15_sp4_h_r_16_46982;
  wire seg_12_15_sp4_h_r_28_43150;
  wire seg_12_15_sp4_h_r_30_43152;
  wire seg_12_15_sp4_h_r_4_50812;
  wire seg_12_15_sp4_r_v_b_3_50451;
  wire seg_12_15_sp4_v_b_17_46746;
  wire seg_12_15_sp4_v_b_20_46749;
  wire seg_12_15_sp4_v_b_31_46870;
  wire seg_12_15_sp4_v_b_6_46625;
  wire seg_12_15_sp4_v_t_38_47112;
  wire seg_12_15_sp4_v_t_43_47117;
  wire seg_12_15_sp4_v_t_46_47120;
  wire seg_12_16_glb_netwk_0_5;
  wire seg_12_16_local_g0_0_50835;
  wire seg_12_16_local_g0_1_50836;
  wire seg_12_16_local_g2_3_50854;
  wire seg_12_16_local_g3_2_50861;
  wire seg_12_16_local_g3_3_50862;
  wire seg_12_16_local_g3_6_50865;
  wire seg_12_16_lutff_1_out_46964;
  wire seg_12_16_lutff_2_out_46965;
  wire seg_12_16_lutff_4_out_46967;
  wire seg_12_16_lutff_5_out_46968;
  wire seg_12_16_lutff_6_out_46969;
  wire seg_12_16_neigh_op_top_1_47087;
  wire seg_12_16_sp4_h_r_16_47105;
  wire seg_12_16_sp4_h_r_8_50939;
  wire seg_12_16_sp4_r_v_b_35_50828;
  wire seg_12_16_sp4_v_b_10_46752;
  wire seg_12_16_sp4_v_b_30_46994;
  wire seg_12_16_sp4_v_b_35_46997;
  wire seg_12_16_sp4_v_b_3_46743;
  wire seg_12_16_sp4_v_b_9_46749;
  wire seg_12_17_glb_netwk_0_5;
  wire seg_12_17_local_g0_2_50960;
  wire seg_12_17_local_g0_4_50962;
  wire seg_12_17_local_g0_5_50963;
  wire seg_12_17_local_g1_1_50967;
  wire seg_12_17_local_g1_5_50971;
  wire seg_12_17_local_g2_6_50980;
  wire seg_12_17_lutff_0_out_47086;
  wire seg_12_17_lutff_1_out_47087;
  wire seg_12_17_lutff_3_out_47089;
  wire seg_12_17_lutff_5_out_47091;
  wire seg_12_17_lutff_6_out_47092;
  wire seg_12_17_neigh_op_bot_4_46967;
  wire seg_12_17_sp4_h_l_39_35732;
  wire seg_12_17_sp4_h_l_41_35734;
  wire seg_12_17_sp4_h_r_10_51054;
  wire seg_12_17_sp4_h_r_1_51053;
  wire seg_12_17_sp4_h_r_21_47231;
  wire seg_12_17_sp4_h_r_2_51056;
  wire seg_12_17_sp4_h_r_38_39564;
  wire seg_12_17_sp4_h_r_7_51061;
  wire seg_12_17_sp4_v_b_10_46875;
  wire seg_12_17_sp4_v_b_5_46868;
  wire seg_12_17_sp4_v_t_37_47357;
  wire seg_12_17_sp4_v_t_41_47361;
  wire seg_12_17_sp4_v_t_44_47364;
  wire seg_12_17_sp4_v_t_45_47365;
  wire seg_12_18_glb_netwk_0_5;
  wire seg_12_18_glb_netwk_1_6;
  wire seg_12_18_local_g0_1_51082;
  wire seg_12_18_local_g0_4_51085;
  wire seg_12_18_local_g0_5_51086;
  wire seg_12_18_local_g0_7_51088;
  wire seg_12_18_local_g1_6_51095;
  wire seg_12_18_local_g2_2_51099;
  wire seg_12_18_local_g2_4_51101;
  wire seg_12_18_local_g2_6_51103;
  wire seg_12_18_local_g3_0_51105;
  wire seg_12_18_local_g3_1_51106;
  wire seg_12_18_lutff_2_out_47211;
  wire seg_12_18_lutff_5_out_47214;
  wire seg_12_18_lutff_7_out_47216;
  wire seg_12_18_neigh_op_lft_4_43382;
  wire seg_12_18_neigh_op_rgt_4_51044;
  wire seg_12_18_neigh_op_top_7_47339;
  wire seg_12_18_sp4_h_l_37_35851;
  wire seg_12_18_sp4_h_l_39_35855;
  wire seg_12_18_sp4_h_l_41_35857;
  wire seg_12_18_sp4_h_l_45_35861;
  wire seg_12_18_sp4_h_l_47_35853;
  wire seg_12_18_sp4_h_r_0_51175;
  wire seg_12_18_sp4_h_r_16_47351;
  wire seg_12_18_sp4_h_r_6_51183;
  wire seg_12_18_sp4_r_v_b_14_50943;
  wire seg_12_18_sp4_r_v_b_16_50945;
  wire seg_12_18_sp4_r_v_b_6_50825;
  wire seg_12_18_sp4_v_b_41_47361;
  wire seg_12_18_sp4_v_b_9_46995;
  wire seg_12_18_sp4_v_t_40_47483;
  wire seg_12_19_glb_netwk_0_5;
  wire seg_12_19_local_g0_6_51210;
  wire seg_12_19_local_g1_1_51213;
  wire seg_12_19_local_g1_2_51214;
  wire seg_12_19_local_g1_3_51215;
  wire seg_12_19_local_g1_4_51216;
  wire seg_12_19_local_g2_0_51220;
  wire seg_12_19_local_g2_2_51222;
  wire seg_12_19_local_g3_0_51228;
  wire seg_12_19_local_g3_3_51231;
  wire seg_12_19_local_g3_7_51235;
  wire seg_12_19_lutff_3_out_47335;
  wire seg_12_19_lutff_4_out_47336;
  wire seg_12_19_lutff_6_out_47338;
  wire seg_12_19_lutff_7_out_47339;
  wire seg_12_19_neigh_op_lft_2_43503;
  wire seg_12_19_neigh_op_top_1_47456;
  wire seg_12_19_sp4_h_l_37_35974;
  wire seg_12_19_sp4_h_l_41_35980;
  wire seg_12_19_sp4_h_l_47_35976;
  wire seg_12_19_sp4_h_r_24_43636;
  wire seg_12_19_sp4_h_r_32_43646;
  wire seg_12_19_sp4_h_r_3_51303;
  wire seg_12_19_sp4_h_r_4_51304;
  wire seg_12_19_sp4_r_v_b_37_51311;
  wire seg_12_19_sp4_v_b_26_47359;
  wire seg_12_19_sp4_v_b_31_47362;
  wire seg_12_19_sp4_v_t_37_47603;
  wire seg_12_20_glb_netwk_0_5;
  wire seg_12_20_glb_netwk_3_8;
  wire seg_12_20_local_g2_0_51343;
  wire seg_12_20_lutff_1_out_47456;
  wire seg_12_20_sp4_v_b_10_47244;
  wire seg_12_20_sp4_v_b_40_47606;
  wire seg_12_20_sp4_v_b_5_47237;
  wire seg_12_21_glb_netwk_0_5;
  wire seg_12_21_local_g0_2_51452;
  wire seg_12_21_local_g0_6_51456;
  wire seg_12_21_local_g1_2_51460;
  wire seg_12_21_local_g1_3_51461;
  wire seg_12_21_local_g2_4_51470;
  wire seg_12_21_local_g2_5_51471;
  wire seg_12_21_local_g2_7_51473;
  wire seg_12_21_local_g3_3_51477;
  wire seg_12_21_lutff_2_out_47580;
  wire seg_12_21_lutff_6_out_47584;
  wire seg_12_21_neigh_op_tnr_3_51535;
  wire seg_12_21_neigh_op_tnr_7_51539;
  wire seg_12_21_sp12_v_b_4_50313;
  wire seg_12_21_sp12_v_t_23_51543;
  wire seg_12_21_sp4_h_r_0_51544;
  wire seg_12_21_sp4_h_r_14_47718;
  wire seg_12_21_sp4_h_r_16_47720;
  wire seg_12_21_sp4_h_r_19_47721;
  wire seg_12_21_sp4_h_r_20_47724;
  wire seg_12_21_sp4_h_r_32_43892;
  wire seg_12_21_sp4_h_r_44_40062;
  wire seg_12_21_sp4_h_r_4_51550;
  wire seg_12_21_sp4_h_r_9_51555;
  wire seg_12_21_sp4_r_v_b_17_51315;
  wire seg_12_21_sp4_r_v_b_1_51187;
  wire seg_12_21_sp4_r_v_b_21_51319;
  wire seg_12_21_sp4_r_v_b_5_51191;
  wire seg_12_21_sp4_r_v_b_9_51195;
  wire seg_12_21_sp4_v_b_0_47357;
  wire seg_12_21_sp4_v_b_10_47367;
  wire seg_12_21_sp4_v_b_16_47483;
  wire seg_12_21_sp4_v_b_1_47356;
  wire seg_12_21_sp4_v_b_37_47726;
  wire seg_12_21_sp4_v_b_4_47361;
  wire seg_12_21_sp4_v_b_8_47365;
  wire seg_12_23_glb_netwk_0_5;
  wire seg_12_23_local_g2_7_51719;
  wire seg_12_23_sp4_h_r_32_44138;
  wire seg_12_23_sp4_h_r_47_40299;
  wire seg_12_23_sp4_r_v_b_1_51433;
  wire seg_12_23_sp4_v_b_0_47603;
  wire seg_12_24_sp4_v_b_6_47732;
  wire seg_12_25_sp4_v_b_1_47848;
  wire seg_12_27_glb_netwk_0_5;
  wire seg_12_27_local_g0_7_52195;
  wire seg_12_27_local_g1_1_52197;
  wire seg_12_27_local_g1_3_52199;
  wire seg_12_27_local_g2_2_52206;
  wire seg_12_27_local_g2_3_52207;
  wire seg_12_27_local_g2_4_52208;
  wire seg_12_27_local_g2_5_52209;
  wire seg_12_27_local_g2_7_52211;
  wire seg_12_27_local_g3_3_52215;
  wire seg_12_27_local_g3_6_52218;
  wire seg_12_27_lutff_2_out_48318;
  wire seg_12_27_lutff_3_out_48319;
  wire seg_12_27_lutff_4_out_48320;
  wire seg_12_27_lutff_5_out_48321;
  wire seg_12_27_lutff_6_out_48322;
  wire seg_12_27_lutff_7_out_48323;
  wire seg_12_27_neigh_op_rgt_4_52151;
  wire seg_12_27_neigh_op_rgt_5_52152;
  wire seg_12_27_neigh_op_rgt_7_52154;
  wire seg_12_27_neigh_op_top_1_48440;
  wire seg_12_27_sp4_h_r_12_48452;
  wire seg_12_27_sp4_h_r_14_48456;
  wire seg_12_27_sp4_r_v_b_19_52055;
  wire seg_12_27_sp4_v_b_19_48224;
  wire seg_12_28_glb_netwk_0_5;
  wire seg_12_28_local_g0_2_52313;
  wire seg_12_28_local_g1_1_52320;
  wire seg_12_28_local_g1_2_52321;
  wire seg_12_28_local_g1_3_52322;
  wire seg_12_28_local_g3_1_52336;
  wire seg_12_28_lutff_1_out_48440;
  wire seg_12_28_lutff_2_out_48441;
  wire seg_12_28_sp4_h_l_43_37089;
  wire seg_12_28_sp4_h_r_10_52407;
  wire seg_12_28_sp4_h_r_11_52408;
  wire seg_12_28_sp4_h_r_18_48583;
  wire seg_12_28_sp4_v_b_9_48225;
  wire seg_12_29_sp4_v_b_1_48340;
  wire seg_12_2_sp4_h_r_6_49215;
  wire seg_12_31_span12_vert_4_51543;
  wire seg_12_31_span4_vert_25_48828;
  wire seg_12_3_sp4_v_t_36_45634;
  wire seg_12_3_sp4_v_t_43_45641;
  wire seg_12_4_sp4_h_l_39_34133;
  wire seg_12_6_sp4_h_l_41_34381;
  wire seg_12_7_sp4_v_t_37_46127;
  wire seg_12_7_sp4_v_t_43_46133;
  wire seg_12_7_sp4_v_t_47_46137;
  wire seg_12_8_glb_netwk_0_5;
  wire seg_12_8_local_g1_3_49862;
  wire seg_12_8_local_g1_7_49866;
  wire seg_12_8_local_g2_5_49872;
  wire seg_12_8_local_g3_0_49875;
  wire seg_12_8_local_g3_1_49876;
  wire seg_12_8_local_g3_5_49880;
  wire seg_12_8_lutff_1_out_45980;
  wire seg_12_8_lutff_5_out_45984;
  wire seg_12_8_neigh_op_bnl_0_42025;
  wire seg_12_8_sp4_h_r_2_49949;
  wire seg_12_8_sp4_h_r_44_38463;
  wire seg_12_8_sp4_r_v_b_31_49840;
  wire seg_12_8_sp4_r_v_b_3_49590;
  wire seg_12_8_sp4_v_b_2_45760;
  wire seg_12_8_sp4_v_b_37_46127;
  wire seg_12_8_sp4_v_b_4_45762;
  wire seg_13_0_local_g1_4_52735;
  wire seg_13_0_local_g1_4_52735_i1;
  wire seg_13_0_local_g1_4_52735_i2;
  wire seg_13_0_local_g1_4_52735_i3;
  wire seg_13_0_span4_horz_r_4_48940;
  wire seg_13_10_sp4_h_l_36_38699;
  wire seg_13_10_sp4_h_l_37_38698;
  wire seg_13_10_sp4_h_r_0_54022;
  wire seg_13_10_sp4_h_r_2_54026;
  wire seg_13_10_sp4_v_b_11_49844;
  wire seg_13_10_sp4_v_t_46_50336;
  wire seg_13_11_glb_netwk_0_5;
  wire seg_13_11_local_g1_5_54064;
  wire seg_13_11_local_g2_2_54069;
  wire seg_13_11_local_g3_6_54081;
  wire seg_13_11_lutff_1_out_50180;
  wire seg_13_11_lutff_6_out_50185;
  wire seg_13_11_sp4_h_l_47_38823;
  wire seg_13_11_sp4_h_r_13_50314;
  wire seg_13_11_sp4_v_b_42_50332;
  wire seg_13_11_sp4_v_t_42_50455;
  wire seg_13_12_glb_netwk_0_5;
  wire seg_13_12_local_g0_1_54175;
  wire seg_13_12_local_g0_2_54176;
  wire seg_13_12_local_g0_3_54177;
  wire seg_13_12_local_g0_4_54178;
  wire seg_13_12_local_g0_5_54179;
  wire seg_13_12_local_g1_4_54186;
  wire seg_13_12_local_g1_5_54187;
  wire seg_13_12_local_g1_6_54188;
  wire seg_13_12_local_g1_7_54189;
  wire seg_13_12_local_g2_0_54190;
  wire seg_13_12_local_g2_1_54191;
  wire seg_13_12_local_g2_3_54193;
  wire seg_13_12_local_g2_5_54195;
  wire seg_13_12_local_g3_4_54202;
  wire seg_13_12_local_g3_7_54205;
  wire seg_13_12_lutff_1_out_50303;
  wire seg_13_12_lutff_2_out_50304;
  wire seg_13_12_lutff_4_out_50306;
  wire seg_13_12_lutff_5_out_50307;
  wire seg_13_12_neigh_op_lft_3_46474;
  wire seg_13_12_neigh_op_lft_4_46475;
  wire seg_13_12_neigh_op_lft_6_46477;
  wire seg_13_12_neigh_op_top_4_50429;
  wire seg_13_12_sp4_h_l_36_38945;
  wire seg_13_12_sp4_h_r_0_54268;
  wire seg_13_12_sp4_h_r_15_50441;
  wire seg_13_12_sp4_h_r_1_54269;
  wire seg_13_12_sp4_h_r_28_46612;
  wire seg_13_12_sp4_h_r_41_42781;
  wire seg_13_12_sp4_h_r_43_42783;
  wire seg_13_12_sp4_h_r_44_42786;
  wire seg_13_12_sp4_h_r_45_42785;
  wire seg_13_12_sp4_h_r_46_42778;
  wire seg_13_12_sp4_h_r_5_54275;
  wire seg_13_12_sp4_h_r_6_54276;
  wire seg_13_12_sp4_r_v_b_23_54045;
  wire seg_13_12_sp4_v_b_10_50091;
  wire seg_13_12_sp4_v_b_18_50209;
  wire seg_13_12_sp4_v_b_21_50212;
  wire seg_13_12_sp4_v_b_24_50327;
  wire seg_13_12_sp4_v_b_9_50088;
  wire seg_13_13_glb_netwk_0_5;
  wire seg_13_13_glb_netwk_1_6;
  wire seg_13_13_local_g0_0_54297;
  wire seg_13_13_local_g0_2_54299;
  wire seg_13_13_local_g0_3_54300;
  wire seg_13_13_local_g0_5_54302;
  wire seg_13_13_local_g1_0_54305;
  wire seg_13_13_local_g1_3_54308;
  wire seg_13_13_local_g1_4_54309;
  wire seg_13_13_local_g1_5_54310;
  wire seg_13_13_local_g1_7_54312;
  wire seg_13_13_local_g2_3_54316;
  wire seg_13_13_local_g2_5_54318;
  wire seg_13_13_local_g2_6_54319;
  wire seg_13_13_local_g3_2_54323;
  wire seg_13_13_local_g3_4_54325;
  wire seg_13_13_local_g3_5_54326;
  wire seg_13_13_local_g3_7_54328;
  wire seg_13_13_lutff_3_out_50428;
  wire seg_13_13_lutff_4_out_50429;
  wire seg_13_13_lutff_5_out_50430;
  wire seg_13_13_lutff_6_out_50431;
  wire seg_13_13_neigh_op_bot_2_50304;
  wire seg_13_13_neigh_op_lft_0_46594;
  wire seg_13_13_neigh_op_lft_3_46597;
  wire seg_13_13_neigh_op_top_4_50552;
  wire seg_13_13_sp4_h_l_37_39067;
  wire seg_13_13_sp4_h_l_45_39077;
  wire seg_13_13_sp4_h_r_0_54391;
  wire seg_13_13_sp4_h_r_16_50567;
  wire seg_13_13_sp4_h_r_23_50562;
  wire seg_13_13_sp4_h_r_2_54395;
  wire seg_13_13_sp4_h_r_30_46737;
  wire seg_13_13_sp4_h_r_37_42898;
  wire seg_13_13_sp4_h_r_43_42906;
  wire seg_13_13_sp4_h_r_44_42909;
  wire seg_13_13_sp4_h_r_46_42901;
  wire seg_13_13_sp4_h_r_4_54397;
  wire seg_13_13_sp4_h_r_5_54398;
  wire seg_13_13_sp4_r_v_b_17_54162;
  wire seg_13_13_sp4_r_v_b_18_54163;
  wire seg_13_13_sp4_r_v_b_23_54168;
  wire seg_13_13_sp4_r_v_b_29_54284;
  wire seg_13_13_sp4_v_b_19_50333;
  wire seg_13_13_sp4_v_t_37_50696;
  wire seg_13_13_sp4_v_t_40_50699;
  wire seg_13_13_sp4_v_t_41_50700;
  wire seg_13_13_sp4_v_t_44_50703;
  wire seg_13_14_glb_netwk_0_5;
  wire seg_13_14_local_g0_6_54426;
  wire seg_13_14_local_g0_7_54427;
  wire seg_13_14_local_g1_0_54428;
  wire seg_13_14_local_g1_3_54431;
  wire seg_13_14_local_g1_5_54433;
  wire seg_13_14_local_g1_6_54434;
  wire seg_13_14_local_g1_7_54435;
  wire seg_13_14_local_g2_1_54437;
  wire seg_13_14_local_g2_6_54442;
  wire seg_13_14_local_g3_0_54444;
  wire seg_13_14_local_g3_2_54446;
  wire seg_13_14_local_g3_3_54447;
  wire seg_13_14_local_g3_5_54449;
  wire seg_13_14_local_g3_6_54450;
  wire seg_13_14_local_g3_7_54451;
  wire seg_13_14_lutff_2_out_50550;
  wire seg_13_14_lutff_3_out_50551;
  wire seg_13_14_lutff_4_out_50552;
  wire seg_13_14_lutff_5_out_50553;
  wire seg_13_14_lutff_7_out_50555;
  wire seg_13_14_neigh_op_bot_5_50430;
  wire seg_13_14_neigh_op_bot_6_50431;
  wire seg_13_14_sp4_h_r_0_54514;
  wire seg_13_14_sp4_h_r_14_50688;
  wire seg_13_14_sp4_h_r_19_50691;
  wire seg_13_14_sp4_h_r_33_46863;
  wire seg_13_14_sp4_h_r_35_46855;
  wire seg_13_14_sp4_r_v_b_13_54281;
  wire seg_13_14_sp4_r_v_b_18_54286;
  wire seg_13_14_sp4_r_v_b_31_54409;
  wire seg_13_14_sp4_r_v_b_3_54159;
  wire seg_13_14_sp4_v_b_0_50327;
  wire seg_13_14_sp4_v_b_23_50460;
  wire seg_13_14_sp4_v_b_30_50579;
  wire seg_13_14_sp4_v_b_38_50697;
  wire seg_13_14_sp4_v_b_40_50699;
  wire seg_13_14_sp4_v_b_6_50333;
  wire seg_13_14_sp4_v_t_40_50822;
  wire seg_13_14_sp4_v_t_41_50823;
  wire seg_13_14_sp4_v_t_42_50824;
  wire seg_13_14_sp4_v_t_44_50826;
  wire seg_13_14_sp4_v_t_45_50827;
  wire seg_13_15_glb_netwk_0_5;
  wire seg_13_15_glb_netwk_3_8;
  wire seg_13_15_local_g0_2_54545;
  wire seg_13_15_local_g0_5_54548;
  wire seg_13_15_local_g1_2_54553;
  wire seg_13_15_local_g1_4_54555;
  wire seg_13_15_local_g2_0_54559;
  wire seg_13_15_local_g2_1_54560;
  wire seg_13_15_local_g2_2_54561;
  wire seg_13_15_local_g2_3_54562;
  wire seg_13_15_local_g2_5_54564;
  wire seg_13_15_local_g2_6_54565;
  wire seg_13_15_local_g3_2_54569;
  wire seg_13_15_local_g3_3_54570;
  wire seg_13_15_local_g3_5_54572;
  wire seg_13_15_local_g3_6_54573;
  wire seg_13_15_lutff_1_out_50672;
  wire seg_13_15_lutff_2_out_50673;
  wire seg_13_15_lutff_4_out_50675;
  wire seg_13_15_lutff_6_out_50677;
  wire seg_13_15_neigh_op_lft_4_46844;
  wire seg_13_15_neigh_op_lft_5_46845;
  wire seg_13_15_neigh_op_rgt_2_54504;
  wire seg_13_15_neigh_op_rgt_6_54508;
  wire seg_13_15_neigh_op_tnl_5_46968;
  wire seg_13_15_neigh_op_tnl_6_46969;
  wire seg_13_15_sp4_h_r_0_54637;
  wire seg_13_15_sp4_h_r_14_50811;
  wire seg_13_15_sp4_h_r_16_50813;
  wire seg_13_15_sp4_h_r_24_46975;
  wire seg_13_15_sp4_h_r_26_46979;
  wire seg_13_15_sp4_h_r_27_46980;
  wire seg_13_15_sp4_h_r_29_46982;
  wire seg_13_15_sp4_h_r_2_54641;
  wire seg_13_15_sp4_r_v_b_23_54414;
  wire seg_13_15_sp4_v_b_26_50698;
  wire seg_13_15_sp4_v_b_43_50825;
  wire seg_13_15_sp4_v_t_41_50946;
  wire seg_13_16_glb_netwk_0_5;
  wire seg_13_16_local_g0_2_54668;
  wire seg_13_16_local_g0_4_54670;
  wire seg_13_16_local_g0_6_54672;
  wire seg_13_16_local_g1_3_54677;
  wire seg_13_16_local_g1_6_54680;
  wire seg_13_16_local_g2_0_54682;
  wire seg_13_16_local_g2_3_54685;
  wire seg_13_16_local_g2_4_54686;
  wire seg_13_16_local_g2_5_54687;
  wire seg_13_16_local_g2_7_54689;
  wire seg_13_16_local_g3_0_54690;
  wire seg_13_16_local_g3_2_54692;
  wire seg_13_16_local_g3_3_54693;
  wire seg_13_16_local_g3_4_54694;
  wire seg_13_16_local_g3_5_54695;
  wire seg_13_16_local_g3_6_54696;
  wire seg_13_16_local_g3_7_54697;
  wire seg_13_16_lutff_1_out_50795;
  wire seg_13_16_neigh_op_bot_4_50675;
  wire seg_13_16_neigh_op_bot_6_50677;
  wire seg_13_16_neigh_op_rgt_0_54625;
  wire seg_13_16_neigh_op_rgt_3_54628;
  wire seg_13_16_neigh_op_rgt_6_54631;
  wire seg_13_16_neigh_op_rgt_7_54632;
  wire seg_13_16_sp4_h_r_11_54763;
  wire seg_13_16_sp4_h_r_22_50932;
  wire seg_13_16_sp4_h_r_24_47098;
  wire seg_13_16_sp4_h_r_26_47102;
  wire seg_13_16_sp4_h_r_27_47103;
  wire seg_13_16_sp4_h_r_2_54764;
  wire seg_13_16_sp4_h_r_31_47107;
  wire seg_13_16_sp4_h_r_34_47100;
  wire seg_13_16_sp4_h_r_37_43267;
  wire seg_13_16_sp4_h_r_44_43278;
  wire seg_13_16_sp4_r_v_b_12_54526;
  wire seg_13_16_sp4_r_v_b_13_54527;
  wire seg_13_16_sp4_r_v_b_21_54535;
  wire seg_13_16_sp4_r_v_b_41_54777;
  wire seg_13_16_sp4_r_v_b_5_54407;
  wire seg_13_16_sp4_r_v_b_7_54409;
  wire seg_13_16_sp4_v_b_0_50573;
  wire seg_13_16_sp4_v_b_14_50697;
  wire seg_13_16_sp4_v_t_43_51071;
  wire seg_13_16_sp4_v_t_46_51074;
  wire seg_13_17_glb_netwk_0_5;
  wire seg_13_17_local_g0_0_54789;
  wire seg_13_17_local_g0_3_54792;
  wire seg_13_17_local_g0_4_54793;
  wire seg_13_17_local_g0_6_54795;
  wire seg_13_17_local_g1_0_54797;
  wire seg_13_17_local_g1_4_54801;
  wire seg_13_17_local_g1_6_54803;
  wire seg_13_17_local_g2_0_54805;
  wire seg_13_17_local_g2_1_54806;
  wire seg_13_17_local_g2_3_54808;
  wire seg_13_17_local_g2_6_54811;
  wire seg_13_17_local_g2_7_54812;
  wire seg_13_17_local_g3_1_54814;
  wire seg_13_17_local_g3_2_54815;
  wire seg_13_17_local_g3_3_54816;
  wire seg_13_17_local_g3_5_54818;
  wire seg_13_17_local_g3_7_54820;
  wire seg_13_17_lutff_6_out_50923;
  wire seg_13_17_neigh_op_bnl_1_46964;
  wire seg_13_17_neigh_op_lft_0_47086;
  wire seg_13_17_neigh_op_lft_3_47089;
  wire seg_13_17_neigh_op_lft_6_47092;
  wire seg_13_17_neigh_op_rgt_2_54750;
  wire seg_13_17_neigh_op_rgt_3_54751;
  wire seg_13_17_neigh_op_rgt_7_54755;
  wire seg_13_17_sp4_h_l_36_39560;
  wire seg_13_17_sp4_h_l_38_39564;
  wire seg_13_17_sp4_h_l_44_39570;
  wire seg_13_17_sp4_h_r_16_51059;
  wire seg_13_17_sp4_h_r_20_51063;
  wire seg_13_17_sp4_h_r_22_51055;
  wire seg_13_17_sp4_h_r_27_47226;
  wire seg_13_17_sp4_h_r_30_47229;
  wire seg_13_17_sp4_h_r_31_47230;
  wire seg_13_17_sp4_h_r_32_47231;
  wire seg_13_17_sp4_h_r_4_54889;
  wire seg_13_17_sp4_h_r_6_54891;
  wire seg_13_17_sp4_r_v_b_11_54536;
  wire seg_13_17_sp4_r_v_b_15_54652;
  wire seg_13_17_sp4_r_v_b_17_54654;
  wire seg_13_17_sp4_r_v_b_21_54658;
  wire seg_13_17_sp4_r_v_b_41_54900;
  wire seg_13_17_sp4_v_b_12_50818;
  wire seg_13_17_sp4_v_b_16_50822;
  wire seg_13_17_sp4_v_b_2_50698;
  wire seg_13_17_sp4_v_t_36_51187;
  wire seg_13_17_sp4_v_t_40_51191;
  wire seg_13_17_sp4_v_t_44_51195;
  wire seg_13_18_glb_netwk_0_5;
  wire seg_13_18_glb_netwk_3_8;
  wire seg_13_18_local_g0_0_54912;
  wire seg_13_18_local_g2_5_54933;
  wire seg_13_18_local_g3_7_54943;
  wire seg_13_18_lutff_3_out_51043;
  wire seg_13_18_lutff_4_out_51044;
  wire seg_13_18_lutff_5_out_51045;
  wire seg_13_18_sp4_h_l_38_39687;
  wire seg_13_18_sp4_h_l_40_39689;
  wire seg_13_18_sp4_h_l_42_39691;
  wire seg_13_18_sp4_h_l_46_39685;
  wire seg_13_18_sp4_r_v_b_13_54773;
  wire seg_13_18_sp4_r_v_b_23_54783;
  wire seg_13_18_sp4_r_v_b_24_54896;
  wire seg_13_18_sp4_v_b_3_50820;
  wire seg_13_18_sp4_v_b_6_50825;
  wire seg_13_18_sp4_v_t_36_51310;
  wire seg_13_18_sp4_v_t_37_51311;
  wire seg_13_18_sp4_v_t_41_51315;
  wire seg_13_18_sp4_v_t_45_51319;
  wire seg_13_19_glb_netwk_0_5;
  wire seg_13_19_glb_netwk_3_8;
  wire seg_13_19_local_g0_7_55042;
  wire seg_13_19_local_g1_0_55043;
  wire seg_13_19_local_g1_6_55049;
  wire seg_13_19_local_g1_7_55050;
  wire seg_13_19_local_g2_1_55052;
  wire seg_13_19_local_g2_2_55053;
  wire seg_13_19_local_g2_4_55055;
  wire seg_13_19_local_g2_5_55056;
  wire seg_13_19_local_g2_6_55057;
  wire seg_13_19_local_g2_7_55058;
  wire seg_13_19_local_g3_3_55062;
  wire seg_13_19_local_g3_4_55063;
  wire seg_13_19_local_g3_5_55064;
  wire seg_13_19_local_g3_7_55066;
  wire seg_13_19_lutff_2_out_51165;
  wire seg_13_19_lutff_6_out_51169;
  wire seg_13_19_lutff_7_out_51170;
  wire seg_13_19_neigh_op_bnl_7_47216;
  wire seg_13_19_neigh_op_rgt_6_55000;
  wire seg_13_19_neigh_op_rgt_7_55001;
  wire seg_13_19_neigh_op_top_0_51286;
  wire seg_13_19_neigh_op_top_7_51293;
  wire seg_13_19_sp4_h_l_36_39806;
  wire seg_13_19_sp4_h_l_38_39810;
  wire seg_13_19_sp4_h_l_40_39812;
  wire seg_13_19_sp4_h_l_41_39811;
  wire seg_13_19_sp4_h_l_44_39816;
  wire seg_13_19_sp4_h_r_18_51307;
  wire seg_13_19_sp4_h_r_2_55133;
  wire seg_13_19_sp4_h_r_41_43642;
  wire seg_13_19_sp4_h_r_8_55139;
  wire seg_13_19_sp4_r_v_b_21_54904;
  wire seg_13_19_sp4_r_v_b_25_55018;
  wire seg_13_19_sp4_v_b_29_51191;
  wire seg_13_19_sp4_v_b_43_51317;
  wire seg_13_19_sp4_v_b_44_51318;
  wire seg_13_19_sp4_v_t_36_51433;
  wire seg_13_20_glb_netwk_0_5;
  wire seg_13_20_local_g1_3_55169;
  wire seg_13_20_local_g1_5_55171;
  wire seg_13_20_local_g1_6_55172;
  wire seg_13_20_local_g2_1_55175;
  wire seg_13_20_local_g2_2_55176;
  wire seg_13_20_local_g2_4_55178;
  wire seg_13_20_local_g2_7_55181;
  wire seg_13_20_local_g3_0_55182;
  wire seg_13_20_local_g3_1_55183;
  wire seg_13_20_local_g3_4_55186;
  wire seg_13_20_local_g3_5_55187;
  wire seg_13_20_local_g3_7_55189;
  wire seg_13_20_lutff_0_out_51286;
  wire seg_13_20_lutff_1_out_51287;
  wire seg_13_20_lutff_4_out_51290;
  wire seg_13_20_lutff_5_out_51291;
  wire seg_13_20_lutff_6_out_51292;
  wire seg_13_20_lutff_7_out_51293;
  wire seg_13_20_neigh_op_tnl_2_47580;
  wire seg_13_20_sp12_v_b_23_55128;
  wire seg_13_20_sp4_h_l_42_39937;
  wire seg_13_20_sp4_h_l_46_39931;
  wire seg_13_20_sp4_h_r_22_51424;
  wire seg_13_20_sp4_h_r_28_47596;
  wire seg_13_20_sp4_h_r_32_47600;
  wire seg_13_20_sp4_h_r_36_43760;
  wire seg_13_20_sp4_h_r_37_43759;
  wire seg_13_20_sp4_h_r_39_43763;
  wire seg_13_20_sp4_h_r_41_43765;
  wire seg_13_20_sp4_h_r_6_55260;
  wire seg_13_20_sp4_v_b_0_51065;
  wire seg_13_20_sp4_v_b_19_51194;
  wire seg_13_20_sp4_v_b_6_51071;
  wire seg_13_21_local_g3_4_55309;
  wire seg_13_21_lutff_6_out_51415;
  wire seg_13_21_sp12_v_b_20_55128;
  wire seg_13_21_sp4_h_r_1_55376;
  wire seg_13_21_sp4_v_b_12_51310;
  wire seg_13_21_sp4_v_b_1_51187;
  wire seg_13_21_sp4_v_t_38_51681;
  wire seg_13_22_glb_netwk_0_5;
  wire seg_13_22_local_g0_1_55405;
  wire seg_13_22_local_g1_5_55417;
  wire seg_13_22_local_g1_6_55418;
  wire seg_13_22_local_g2_2_55422;
  wire seg_13_22_local_g2_3_55423;
  wire seg_13_22_local_g3_5_55433;
  wire seg_13_22_lutff_1_out_51533;
  wire seg_13_22_lutff_3_out_51535;
  wire seg_13_22_lutff_5_out_51537;
  wire seg_13_22_lutff_7_out_51539;
  wire seg_13_22_neigh_op_bot_6_51415;
  wire seg_13_22_sp12_v_b_19_55128;
  wire seg_13_22_sp12_v_b_21_55250;
  wire seg_13_22_sp4_h_r_26_47840;
  wire seg_13_22_sp4_v_b_38_51681;
  wire seg_13_24_sp4_v_b_8_51565;
  wire seg_13_27_glb_netwk_0_5;
  wire seg_13_27_local_g0_2_56021;
  wire seg_13_27_local_g0_5_56024;
  wire seg_13_27_local_g0_6_56025;
  wire seg_13_27_local_g0_7_56026;
  wire seg_13_27_local_g1_3_56030;
  wire seg_13_27_local_g1_4_56031;
  wire seg_13_27_local_g1_7_56034;
  wire seg_13_27_local_g2_1_56036;
  wire seg_13_27_local_g2_2_56037;
  wire seg_13_27_local_g2_5_56040;
  wire seg_13_27_local_g3_4_56047;
  wire seg_13_27_lutff_2_out_52149;
  wire seg_13_27_lutff_4_out_52151;
  wire seg_13_27_lutff_5_out_52152;
  wire seg_13_27_lutff_7_out_52154;
  wire seg_13_27_neigh_op_lft_4_48320;
  wire seg_13_27_neigh_op_lft_5_48321;
  wire seg_13_27_neigh_op_lft_6_48322;
  wire seg_13_27_neigh_op_lft_7_48323;
  wire seg_13_27_neigh_op_tnl_1_48440;
  wire seg_13_27_sp4_r_v_b_13_55880;
  wire seg_13_27_sp4_v_b_18_52054;
  wire seg_13_27_sp4_v_b_19_52055;
  wire seg_13_28_sp4_h_r_6_56244;
  wire seg_13_28_sp4_h_r_7_56245;
  wire seg_13_28_sp4_v_b_4_52053;
  wire seg_13_2_sp4_h_l_46_37717;
  wire seg_13_31_glb_netwk_0_5;
  wire seg_13_31_local_g1_2_56534;
  wire seg_13_31_local_g1_3_56535;
  wire seg_13_31_local_g1_4_56536;
  wire seg_13_31_local_g1_4_56536_i1;
  wire seg_13_31_local_g1_4_56536_i2;
  wire seg_13_31_local_g1_4_56536_i3;
  wire seg_13_31_span12_vert_0_55128;
  wire seg_13_31_span12_vert_2_55250;
  wire seg_13_31_span4_horz_r_11_48881;
  wire seg_13_31_span4_horz_r_4_52709;
  wire seg_13_31_span4_vert_18_52546;
  wire seg_13_3_glb_netwk_0_5;
  wire seg_13_3_local_g0_6_53073;
  wire seg_13_3_local_g0_7_53074;
  wire seg_13_3_local_g1_3_53078;
  wire seg_13_3_local_g3_1_53092;
  wire seg_13_3_local_g3_4_53095;
  wire seg_13_3_local_g3_7_53098;
  wire seg_13_3_lutff_7_out_49202;
  wire seg_13_3_neigh_op_tnr_1_53150;
  wire seg_13_3_neigh_op_tnr_4_53153;
  wire seg_13_3_neigh_op_top_6_49324;
  wire seg_13_3_neigh_op_top_7_49325;
  wire seg_13_3_sp4_h_r_11_53164;
  wire seg_13_3_sp4_r_v_b_19_52929;
  wire seg_13_3_sp4_r_v_b_23_52933;
  wire seg_13_3_sp4_v_t_43_49472;
  wire seg_13_3_sp4_v_t_46_49475;
  wire seg_13_4_glb_netwk_0_5;
  wire seg_13_4_local_g0_4_53194;
  wire seg_13_4_local_g1_0_53198;
  wire seg_13_4_local_g1_6_53204;
  wire seg_13_4_local_g2_2_53208;
  wire seg_13_4_local_g2_4_53210;
  wire seg_13_4_local_g2_5_53211;
  wire seg_13_4_local_g2_7_53213;
  wire seg_13_4_local_g3_0_53214;
  wire seg_13_4_local_g3_1_53215;
  wire seg_13_4_local_g3_7_53221;
  wire seg_13_4_lutff_2_out_49320;
  wire seg_13_4_lutff_3_out_49321;
  wire seg_13_4_lutff_4_out_49322;
  wire seg_13_4_lutff_5_out_49323;
  wire seg_13_4_lutff_6_out_49324;
  wire seg_13_4_lutff_7_out_49325;
  wire seg_13_4_neigh_op_bnr_0_53026;
  wire seg_13_4_neigh_op_rgt_0_53149;
  wire seg_13_4_neigh_op_rgt_1_53150;
  wire seg_13_4_neigh_op_rgt_2_53151;
  wire seg_13_4_neigh_op_rgt_4_53153;
  wire seg_13_4_neigh_op_rgt_7_53156;
  wire seg_13_4_sp4_h_l_44_37971;
  wire seg_13_6_sp4_h_l_46_38209;
  wire seg_13_7_sp4_v_t_38_49959;
  wire seg_13_8_local_g0_0_53682;
  wire seg_13_8_local_g0_1_53683;
  wire seg_13_8_local_g0_5_53687;
  wire seg_13_8_local_g0_6_53688;
  wire seg_13_8_local_g1_0_53690;
  wire seg_13_8_local_g1_6_53696;
  wire seg_13_8_local_g3_6_53712;
  wire seg_13_8_local_g3_7_53713;
  wire seg_13_8_lutff_2_out_49812;
  wire seg_13_8_lutff_3_out_49813;
  wire seg_13_8_lutff_4_out_49814;
  wire seg_13_8_lutff_5_out_49815;
  wire seg_13_8_lutff_7_out_49817;
  wire seg_13_8_neigh_op_bnr_6_53524;
  wire seg_13_8_neigh_op_rgt_6_53647;
  wire seg_13_8_neigh_op_rgt_7_53648;
  wire seg_13_8_neigh_op_top_0_49933;
  wire seg_13_8_neigh_op_top_1_49934;
  wire seg_13_8_neigh_op_top_5_49938;
  wire seg_13_8_neigh_op_top_6_49939;
  wire seg_13_8_sp4_h_l_44_38463;
  wire seg_13_8_sp4_h_r_12_49946;
  wire seg_13_8_sp4_h_r_8_53786;
  wire seg_13_8_sp4_v_b_9_49596;
  wire seg_13_9_glb_netwk_0_5;
  wire seg_13_9_local_g0_2_53807;
  wire seg_13_9_local_g0_4_53809;
  wire seg_13_9_local_g1_1_53814;
  wire seg_13_9_local_g1_2_53815;
  wire seg_13_9_local_g1_4_53817;
  wire seg_13_9_local_g1_5_53818;
  wire seg_13_9_local_g1_6_53819;
  wire seg_13_9_local_g1_7_53820;
  wire seg_13_9_local_g2_2_53823;
  wire seg_13_9_local_g2_4_53825;
  wire seg_13_9_local_g2_6_53827;
  wire seg_13_9_local_g3_2_53831;
  wire seg_13_9_local_g3_3_53832;
  wire seg_13_9_local_g3_5_53834;
  wire seg_13_9_local_g3_7_53836;
  wire seg_13_9_lutff_0_out_49933;
  wire seg_13_9_lutff_1_out_49934;
  wire seg_13_9_lutff_5_out_49938;
  wire seg_13_9_lutff_6_out_49939;
  wire seg_13_9_neigh_op_bnr_6_53647;
  wire seg_13_9_neigh_op_bot_2_49812;
  wire seg_13_9_neigh_op_bot_4_49814;
  wire seg_13_9_neigh_op_bot_5_49815;
  wire seg_13_9_neigh_op_bot_7_49817;
  wire seg_13_9_neigh_op_rgt_2_53766;
  wire seg_13_9_neigh_op_rgt_4_53768;
  wire seg_13_9_neigh_op_rgt_5_53769;
  wire seg_13_9_neigh_op_rgt_7_53771;
  wire seg_13_9_sp4_h_r_20_50079;
  wire seg_13_9_sp4_h_r_27_46242;
  wire seg_13_9_sp4_r_v_b_18_53671;
  wire seg_13_9_sp4_r_v_b_21_53674;
  wire seg_13_9_sp4_v_b_18_49840;
  wire seg_14_10_local_g0_5_57763;
  wire seg_14_10_local_g0_6_57764;
  wire seg_14_10_local_g2_2_57776;
  wire seg_14_10_local_g2_5_57779;
  wire seg_14_10_neigh_op_bnr_5_57599;
  wire seg_14_10_sp4_h_l_36_42530;
  wire seg_14_10_sp4_h_l_38_42534;
  wire seg_14_10_sp4_h_l_39_42533;
  wire seg_14_10_sp4_h_r_22_54025;
  wire seg_14_10_sp4_h_r_45_46370;
  wire seg_14_10_sp4_h_r_46_46363;
  wire seg_14_10_sp4_r_v_b_10_57506;
  wire seg_14_10_sp4_v_b_8_53674;
  wire seg_14_11_glb_netwk_0_5;
  wire seg_14_11_glb_netwk_3_8;
  wire seg_14_11_local_g0_3_57884;
  wire seg_14_11_local_g0_4_57885;
  wire seg_14_11_local_g0_6_57887;
  wire seg_14_11_local_g0_7_57888;
  wire seg_14_11_local_g1_1_57890;
  wire seg_14_11_local_g1_4_57893;
  wire seg_14_11_local_g2_0_57897;
  wire seg_14_11_local_g2_2_57899;
  wire seg_14_11_local_g2_3_57900;
  wire seg_14_11_local_g2_5_57902;
  wire seg_14_11_local_g2_6_57903;
  wire seg_14_11_lutff_0_out_54010;
  wire seg_14_11_lutff_1_out_54011;
  wire seg_14_11_lutff_3_out_54013;
  wire seg_14_11_lutff_5_out_54015;
  wire seg_14_11_lutff_6_out_54016;
  wire seg_14_11_lutff_7_out_54017;
  wire seg_14_11_neigh_op_bnr_4_57721;
  wire seg_14_11_neigh_op_lft_6_50185;
  wire seg_14_11_sp12_h_r_4_50310;
  wire seg_14_11_sp4_h_r_11_57978;
  wire seg_14_11_sp4_h_r_24_50314;
  wire seg_14_11_sp4_h_r_26_50318;
  wire seg_14_11_sp4_h_r_4_57981;
  wire seg_14_11_sp4_r_v_b_35_57874;
  wire seg_14_11_sp4_r_v_b_37_57988;
  wire seg_14_11_sp4_v_b_30_54041;
  wire seg_14_11_sp4_v_b_40_54161;
  wire seg_14_11_sp4_v_b_45_54166;
  wire seg_14_11_sp4_v_t_45_54289;
  wire seg_14_12_glb_netwk_0_5;
  wire seg_14_12_local_g0_2_58006;
  wire seg_14_12_local_g0_3_58007;
  wire seg_14_12_local_g1_0_58012;
  wire seg_14_12_local_g1_1_58013;
  wire seg_14_12_local_g1_2_58014;
  wire seg_14_12_local_g1_3_58015;
  wire seg_14_12_local_g1_6_58018;
  wire seg_14_12_local_g1_7_58019;
  wire seg_14_12_local_g2_1_58021;
  wire seg_14_12_local_g2_3_58023;
  wire seg_14_12_local_g2_4_58024;
  wire seg_14_12_local_g2_6_58026;
  wire seg_14_12_local_g2_7_58027;
  wire seg_14_12_local_g3_3_58031;
  wire seg_14_12_local_g3_6_58034;
  wire seg_14_12_local_g3_7_58035;
  wire seg_14_12_lutff_1_out_54134;
  wire seg_14_12_lutff_2_out_54135;
  wire seg_14_12_lutff_3_out_54136;
  wire seg_14_12_lutff_6_out_54139;
  wire seg_14_12_neigh_op_bnr_1_57841;
  wire seg_14_12_neigh_op_bnr_2_57842;
  wire seg_14_12_neigh_op_bnr_7_57847;
  wire seg_14_12_neigh_op_bot_3_54013;
  wire seg_14_12_sp4_h_l_38_42780;
  wire seg_14_12_sp4_h_r_28_50443;
  wire seg_14_12_sp4_h_r_2_58102;
  wire seg_14_12_sp4_h_r_39_46610;
  wire seg_14_12_sp4_h_r_40_46613;
  wire seg_14_12_sp4_h_r_42_46615;
  wire seg_14_12_sp4_h_r_43_46614;
  wire seg_14_12_sp4_r_v_b_0_57742;
  wire seg_14_12_sp4_r_v_b_14_57866;
  wire seg_14_12_sp4_r_v_b_15_57867;
  wire seg_14_12_sp4_r_v_b_30_57994;
  wire seg_14_12_sp4_r_v_b_31_57993;
  wire seg_14_12_sp4_r_v_b_33_57995;
  wire seg_14_12_sp4_v_b_18_54040;
  wire seg_14_12_sp4_v_b_19_54041;
  wire seg_14_12_sp4_v_b_27_54159;
  wire seg_14_12_sp4_v_b_39_54283;
  wire seg_14_12_sp4_v_b_4_53916;
  wire seg_14_13_glb_netwk_0_5;
  wire seg_14_13_local_g0_1_58128;
  wire seg_14_13_local_g0_2_58129;
  wire seg_14_13_local_g0_3_58130;
  wire seg_14_13_local_g0_6_58133;
  wire seg_14_13_local_g0_7_58134;
  wire seg_14_13_local_g1_0_58135;
  wire seg_14_13_local_g1_1_58136;
  wire seg_14_13_local_g1_2_58137;
  wire seg_14_13_local_g1_3_58138;
  wire seg_14_13_local_g1_5_58140;
  wire seg_14_13_local_g1_6_58141;
  wire seg_14_13_local_g1_7_58142;
  wire seg_14_13_local_g2_1_58144;
  wire seg_14_13_local_g2_2_58145;
  wire seg_14_13_local_g2_4_58147;
  wire seg_14_13_local_g2_5_58148;
  wire seg_14_13_local_g2_6_58149;
  wire seg_14_13_local_g2_7_58150;
  wire seg_14_13_local_g3_0_58151;
  wire seg_14_13_local_g3_1_58152;
  wire seg_14_13_local_g3_3_58154;
  wire seg_14_13_local_g3_4_58155;
  wire seg_14_13_local_g3_5_58156;
  wire seg_14_13_local_g3_6_58157;
  wire seg_14_13_local_g3_7_58158;
  wire seg_14_13_lutff_2_out_54258;
  wire seg_14_13_lutff_7_out_54263;
  wire seg_14_13_neigh_op_bnl_1_50303;
  wire seg_14_13_neigh_op_bnr_1_57964;
  wire seg_14_13_neigh_op_bnr_6_57969;
  wire seg_14_13_neigh_op_bnr_7_57970;
  wire seg_14_13_neigh_op_bot_2_54135;
  wire seg_14_13_neigh_op_bot_3_54136;
  wire seg_14_13_neigh_op_lft_3_50428;
  wire seg_14_13_sp12_h_r_9_42895;
  wire seg_14_13_sp4_h_l_36_42899;
  wire seg_14_13_sp4_h_l_41_42904;
  wire seg_14_13_sp4_h_r_10_58223;
  wire seg_14_13_sp4_h_r_16_54398;
  wire seg_14_13_sp4_h_r_24_50560;
  wire seg_14_13_sp4_h_r_26_50564;
  wire seg_14_13_sp4_h_r_27_50565;
  wire seg_14_13_sp4_h_r_2_58225;
  wire seg_14_13_sp4_h_r_30_50568;
  wire seg_14_13_sp4_h_r_32_50570;
  wire seg_14_13_sp4_h_r_39_46733;
  wire seg_14_13_sp4_h_r_41_46735;
  wire seg_14_13_sp4_h_r_6_58229;
  wire seg_14_13_sp4_h_r_8_58231;
  wire seg_14_13_sp4_r_v_b_12_57987;
  wire seg_14_13_sp4_r_v_b_21_57996;
  wire seg_14_13_sp4_r_v_b_26_58113;
  wire seg_14_13_sp4_r_v_b_30_58117;
  wire seg_14_13_sp4_r_v_b_39_58236;
  wire seg_14_13_sp4_r_v_b_5_57868;
  wire seg_14_13_sp4_v_b_12_54157;
  wire seg_14_13_sp4_v_b_28_54285;
  wire seg_14_13_sp4_v_b_34_54291;
  wire seg_14_13_sp4_v_b_38_54405;
  wire seg_14_13_sp4_v_b_40_54407;
  wire seg_14_13_sp4_v_b_45_54412;
  wire seg_14_13_sp4_v_b_47_54414;
  wire seg_14_13_sp4_v_t_37_54527;
  wire seg_14_13_sp4_v_t_41_54531;
  wire seg_14_13_sp4_v_t_43_54533;
  wire seg_14_14_glb_netwk_0_5;
  wire seg_14_14_glb_netwk_3_8;
  wire seg_14_14_local_g1_0_58258;
  wire seg_14_14_local_g1_2_58260;
  wire seg_14_14_local_g1_3_58261;
  wire seg_14_14_local_g1_4_58262;
  wire seg_14_14_local_g1_5_58263;
  wire seg_14_14_local_g1_6_58264;
  wire seg_14_14_local_g2_4_58270;
  wire seg_14_14_local_g2_6_58272;
  wire seg_14_14_local_g2_7_58273;
  wire seg_14_14_local_g3_0_58274;
  wire seg_14_14_local_g3_2_58276;
  wire seg_14_14_local_g3_3_58277;
  wire seg_14_14_local_g3_5_58279;
  wire seg_14_14_local_g3_6_58280;
  wire seg_14_14_local_g3_7_58281;
  wire seg_14_14_lutff_1_out_54380;
  wire seg_14_14_lutff_5_out_54384;
  wire seg_14_14_lutff_6_out_54385;
  wire seg_14_14_neigh_op_lft_3_50551;
  wire seg_14_14_neigh_op_top_0_54502;
  wire seg_14_14_neigh_op_top_4_54506;
  wire seg_14_14_sp4_h_l_36_43022;
  wire seg_14_14_sp4_h_l_38_43026;
  wire seg_14_14_sp4_h_l_40_43028;
  wire seg_14_14_sp4_h_l_47_43023;
  wire seg_14_14_sp4_h_r_0_58344;
  wire seg_14_14_sp4_h_r_14_54519;
  wire seg_14_14_sp4_h_r_20_54525;
  wire seg_14_14_sp4_h_r_39_46856;
  wire seg_14_14_sp4_h_r_40_46859;
  wire seg_14_14_sp4_h_r_44_46863;
  wire seg_14_14_sp4_h_r_6_58352;
  wire seg_14_14_sp4_r_v_b_19_58117;
  wire seg_14_14_sp4_r_v_b_23_58121;
  wire seg_14_14_sp4_r_v_b_2_57990;
  wire seg_14_14_sp4_r_v_b_33_58241;
  wire seg_14_14_sp4_v_b_14_54282;
  wire seg_14_14_sp4_v_b_1_54157;
  wire seg_14_14_sp4_v_b_20_54288;
  wire seg_14_14_sp4_v_b_26_54406;
  wire seg_14_14_sp4_v_b_46_54536;
  wire seg_14_14_sp4_v_b_47_54537;
  wire seg_14_14_sp4_v_b_4_54162;
  wire seg_14_14_sp4_v_b_5_54161;
  wire seg_14_14_sp4_v_b_8_54166;
  wire seg_14_15_glb_netwk_0_5;
  wire seg_14_15_local_g1_1_58382;
  wire seg_14_15_local_g1_2_58383;
  wire seg_14_15_local_g1_5_58386;
  wire seg_14_15_local_g1_6_58387;
  wire seg_14_15_local_g2_2_58391;
  wire seg_14_15_local_g2_3_58392;
  wire seg_14_15_local_g2_6_58395;
  wire seg_14_15_local_g2_7_58396;
  wire seg_14_15_local_g3_0_58397;
  wire seg_14_15_local_g3_1_58398;
  wire seg_14_15_local_g3_5_58402;
  wire seg_14_15_local_g3_6_58403;
  wire seg_14_15_local_g3_7_58404;
  wire seg_14_15_lutff_0_out_54502;
  wire seg_14_15_lutff_2_out_54504;
  wire seg_14_15_lutff_4_out_54506;
  wire seg_14_15_lutff_6_out_54508;
  wire seg_14_15_lutff_7_out_54509;
  wire seg_14_15_neigh_op_tnl_1_50795;
  wire seg_14_15_sp4_h_r_14_54642;
  wire seg_14_15_sp4_h_r_30_50814;
  wire seg_14_15_sp4_h_r_35_50809;
  wire seg_14_15_sp4_h_r_45_46985;
  wire seg_14_15_sp4_h_r_47_46977;
  wire seg_14_15_sp4_r_v_b_16_58237;
  wire seg_14_15_sp4_r_v_b_23_58244;
  wire seg_14_15_sp4_r_v_b_25_58356;
  wire seg_14_15_sp4_r_v_b_29_58360;
  wire seg_14_15_sp4_r_v_b_2_58113;
  wire seg_14_15_sp4_v_b_0_54281;
  wire seg_14_15_sp4_v_b_10_54291;
  wire seg_14_15_sp4_v_b_26_54529;
  wire seg_14_15_sp4_v_b_2_54283;
  wire seg_14_15_sp4_v_b_30_54533;
  wire seg_14_15_sp4_v_b_39_54652;
  wire seg_14_15_sp4_v_b_3_54282;
  wire seg_14_15_sp4_v_b_4_54285;
  wire seg_14_15_sp4_v_b_9_54288;
  wire seg_14_15_sp4_v_t_40_54776;
  wire seg_14_15_sp4_v_t_41_54777;
  wire seg_14_15_sp4_v_t_46_54782;
  wire seg_14_16_glb_netwk_0_5;
  wire seg_14_16_local_g0_2_58498;
  wire seg_14_16_local_g0_4_58500;
  wire seg_14_16_local_g0_5_58501;
  wire seg_14_16_local_g1_0_58504;
  wire seg_14_16_local_g1_5_58509;
  wire seg_14_16_local_g1_7_58511;
  wire seg_14_16_local_g2_1_58513;
  wire seg_14_16_local_g2_5_58517;
  wire seg_14_16_local_g2_6_58518;
  wire seg_14_16_local_g3_0_58520;
  wire seg_14_16_local_g3_1_58521;
  wire seg_14_16_local_g3_3_58523;
  wire seg_14_16_lutff_0_out_54625;
  wire seg_14_16_lutff_3_out_54628;
  wire seg_14_16_lutff_5_out_54630;
  wire seg_14_16_lutff_6_out_54631;
  wire seg_14_16_lutff_7_out_54632;
  wire seg_14_16_neigh_op_bot_0_54502;
  wire seg_14_16_neigh_op_bot_4_54506;
  wire seg_14_16_neigh_op_bot_7_54509;
  wire seg_14_16_neigh_op_tnl_6_50923;
  wire seg_14_16_sp4_h_r_25_50930;
  wire seg_14_16_sp4_h_r_32_50939;
  wire seg_14_16_sp4_h_r_41_47104;
  wire seg_14_16_sp4_r_v_b_13_58357;
  wire seg_14_16_sp4_r_v_b_33_58487;
  wire seg_14_16_sp4_r_v_b_43_58609;
  wire seg_14_16_sp4_r_v_b_5_58237;
  wire seg_14_16_sp4_v_b_0_54404;
  wire seg_14_16_sp4_v_b_2_54406;
  wire seg_14_16_sp4_v_b_8_54412;
  wire seg_14_16_sp4_v_t_41_54900;
  wire seg_14_17_glb_netwk_0_5;
  wire seg_14_17_local_g0_1_58620;
  wire seg_14_17_local_g1_3_58630;
  wire seg_14_17_local_g1_6_58633;
  wire seg_14_17_local_g3_1_58644;
  wire seg_14_17_local_g3_2_58645;
  wire seg_14_17_local_g3_7_58650;
  wire seg_14_17_lutff_1_out_54749;
  wire seg_14_17_lutff_2_out_54750;
  wire seg_14_17_lutff_3_out_54751;
  wire seg_14_17_lutff_7_out_54755;
  wire seg_14_17_neigh_op_rgt_2_58580;
  wire seg_14_17_neigh_op_rgt_7_58585;
  wire seg_14_17_sp4_h_l_42_43399;
  wire seg_14_17_sp4_h_l_43_43398;
  wire seg_14_17_sp4_h_l_45_43400;
  wire seg_14_17_sp4_h_r_11_58716;
  wire seg_14_17_sp4_r_v_b_30_58609;
  wire seg_14_17_sp4_v_b_10_54537;
  wire seg_14_17_sp4_v_b_17_54654;
  wire seg_14_17_sp4_v_t_36_55018;
  wire seg_14_17_sp4_v_t_43_55025;
  wire seg_14_17_sp4_v_t_45_55027;
  wire seg_14_18_glb_netwk_0_5;
  wire seg_14_18_local_g0_3_58745;
  wire seg_14_18_local_g0_5_58747;
  wire seg_14_18_local_g0_7_58749;
  wire seg_14_18_local_g1_3_58753;
  wire seg_14_18_local_g2_0_58758;
  wire seg_14_18_local_g2_1_58759;
  wire seg_14_18_local_g2_2_58760;
  wire seg_14_18_local_g2_3_58761;
  wire seg_14_18_local_g2_5_58763;
  wire seg_14_18_local_g2_6_58764;
  wire seg_14_18_local_g3_0_58766;
  wire seg_14_18_local_g3_1_58767;
  wire seg_14_18_local_g3_3_58769;
  wire seg_14_18_lutff_0_out_54871;
  wire seg_14_18_lutff_1_out_54872;
  wire seg_14_18_lutff_3_out_54874;
  wire seg_14_18_lutff_5_out_54876;
  wire seg_14_18_neigh_op_lft_3_51043;
  wire seg_14_18_neigh_op_lft_5_51045;
  wire seg_14_18_neigh_op_tnr_3_58827;
  wire seg_14_18_sp4_h_l_41_43519;
  wire seg_14_18_sp4_h_l_45_43523;
  wire seg_14_18_sp4_h_r_14_55011;
  wire seg_14_18_sp4_h_r_41_47350;
  wire seg_14_18_sp4_h_r_8_58846;
  wire seg_14_18_sp4_h_r_9_58847;
  wire seg_14_18_sp4_r_v_b_10_58490;
  wire seg_14_18_sp4_r_v_b_41_58853;
  wire seg_14_18_sp4_v_b_10_54660;
  wire seg_14_18_sp4_v_b_23_54783;
  wire seg_14_18_sp4_v_b_24_54896;
  wire seg_14_18_sp4_v_b_38_55020;
  wire seg_14_18_sp4_v_b_43_55025;
  wire seg_14_19_glb_netwk_0_5;
  wire seg_14_19_glb_netwk_1_6;
  wire seg_14_19_local_g0_0_58865;
  wire seg_14_19_local_g0_2_58867;
  wire seg_14_19_local_g1_0_58873;
  wire seg_14_19_local_g1_2_58875;
  wire seg_14_19_local_g1_4_58877;
  wire seg_14_19_local_g2_3_58884;
  wire seg_14_19_local_g3_3_58892;
  wire seg_14_19_local_g3_5_58894;
  wire seg_14_19_lutff_0_out_54994;
  wire seg_14_19_lutff_1_out_54995;
  wire seg_14_19_lutff_6_out_55000;
  wire seg_14_19_lutff_7_out_55001;
  wire seg_14_19_neigh_op_rgt_3_58827;
  wire seg_14_19_neigh_op_top_0_55117;
  wire seg_14_19_neigh_op_top_4_55121;
  wire seg_14_19_sp4_h_l_37_43636;
  wire seg_14_19_sp4_h_l_39_43640;
  wire seg_14_19_sp4_h_l_43_43644;
  wire seg_14_19_sp4_h_l_47_43638;
  wire seg_14_19_sp4_h_r_10_58961;
  wire seg_14_19_sp4_h_r_11_58962;
  wire seg_14_19_sp4_h_r_43_47475;
  wire seg_14_19_sp4_r_v_b_21_58734;
  wire seg_14_19_sp4_r_v_b_33_58856;
  wire seg_14_19_sp4_v_t_39_55267;
  wire seg_14_20_glb_netwk_0_5;
  wire seg_14_20_local_g0_0_58988;
  wire seg_14_20_local_g0_2_58990;
  wire seg_14_20_local_g0_3_58991;
  wire seg_14_20_local_g0_4_58992;
  wire seg_14_20_local_g0_5_58993;
  wire seg_14_20_local_g0_6_58994;
  wire seg_14_20_local_g0_7_58995;
  wire seg_14_20_local_g1_3_58999;
  wire seg_14_20_local_g1_6_59002;
  wire seg_14_20_local_g2_0_59004;
  wire seg_14_20_local_g2_1_59005;
  wire seg_14_20_local_g3_2_59014;
  wire seg_14_20_local_g3_4_59016;
  wire seg_14_20_local_g3_5_59017;
  wire seg_14_20_lutff_0_out_55117;
  wire seg_14_20_lutff_1_out_55118;
  wire seg_14_20_lutff_2_out_55119;
  wire seg_14_20_lutff_4_out_55121;
  wire seg_14_20_neigh_op_bnr_3_58827;
  wire seg_14_20_neigh_op_lft_4_51290;
  wire seg_14_20_neigh_op_lft_6_51292;
  wire seg_14_20_neigh_op_top_7_55247;
  wire seg_14_20_sp4_h_l_37_43759;
  wire seg_14_20_sp4_h_l_39_43763;
  wire seg_14_20_sp4_h_l_41_43765;
  wire seg_14_20_sp4_h_l_43_43767;
  wire seg_14_20_sp4_h_r_0_59082;
  wire seg_14_20_sp4_h_r_10_59084;
  wire seg_14_20_sp4_h_r_18_55261;
  wire seg_14_20_sp4_h_r_45_47600;
  wire seg_14_20_sp4_h_r_5_59089;
  wire seg_14_20_sp4_r_v_b_20_58856;
  wire seg_14_20_sp4_r_v_b_27_58973;
  wire seg_14_20_sp4_r_v_b_6_58732;
  wire seg_14_20_sp4_r_v_b_8_58734;
  wire seg_14_20_sp4_v_b_14_55020;
  wire seg_14_20_sp4_v_b_19_55025;
  wire seg_14_20_sp4_v_b_3_54897;
  wire seg_14_21_glb_netwk_0_5;
  wire seg_14_21_glb_netwk_1_6;
  wire seg_14_21_local_g3_5_59140;
  wire seg_14_21_lutff_7_out_55247;
  wire seg_14_21_sp4_h_l_45_43892;
  wire seg_14_21_sp4_h_r_1_59206;
  wire seg_14_21_sp4_v_b_37_55388;
  wire seg_14_22_sp4_v_b_3_55143;
  wire seg_14_22_sp4_v_b_6_55148;
  wire seg_14_23_sp4_h_l_45_44138;
  wire seg_14_24_sp4_v_b_11_55397;
  wire seg_14_25_sp4_h_r_9_59708;
  wire seg_14_26_glb_netwk_0_5;
  wire seg_14_26_local_g1_1_59735;
  wire seg_14_26_local_g1_3_59737;
  wire seg_14_26_local_g3_3_59753;
  wire seg_14_26_lutff_3_out_55858;
  wire seg_14_26_sp4_r_v_b_25_59709;
  wire seg_14_26_sp4_v_b_11_55643;
  wire seg_14_26_sp4_v_b_9_55641;
  wire seg_14_27_glb_netwk_0_5;
  wire seg_14_27_local_g0_2_59851;
  wire seg_14_27_local_g1_2_59859;
  wire seg_14_27_local_g1_5_59862;
  wire seg_14_27_local_g2_2_59867;
  wire seg_14_27_local_g2_4_59869;
  wire seg_14_27_local_g2_5_59870;
  wire seg_14_27_local_g3_2_59875;
  wire seg_14_27_local_g3_6_59879;
  wire seg_14_27_lutff_2_out_55980;
  wire seg_14_27_lutff_5_out_55983;
  wire seg_14_27_neigh_op_lft_5_52152;
  wire seg_14_27_sp4_h_r_36_48452;
  wire seg_14_27_sp4_h_r_38_48456;
  wire seg_14_27_sp4_r_v_b_10_59597;
  wire seg_14_27_sp4_r_v_b_18_59715;
  wire seg_14_27_sp4_r_v_b_35_59842;
  wire seg_14_27_sp4_v_b_18_55885;
  wire seg_14_28_local_g1_4_59984;
  wire seg_14_28_local_g2_0_59988;
  wire seg_14_28_neigh_op_rgt_0_59931;
  wire seg_14_28_sp4_h_r_18_56245;
  wire seg_14_28_sp4_h_r_34_52407;
  wire seg_14_28_sp4_v_b_0_55880;
  wire seg_14_28_sp4_v_b_20_56010;
  wire seg_14_2_local_g0_2_56776;
  wire seg_14_2_local_g0_3_56777;
  wire seg_14_2_local_g0_6_56780;
  wire seg_14_2_local_g1_3_56785;
  wire seg_14_2_local_g2_0_56790;
  wire seg_14_2_local_g2_3_56793;
  wire seg_14_2_local_g3_2_56800;
  wire seg_14_2_local_g3_7_56805;
  wire seg_14_2_lutff_2_out_52869;
  wire seg_14_2_lutff_3_out_52870;
  wire seg_14_2_neigh_op_rgt_0_56697;
  wire seg_14_2_neigh_op_tnr_2_56858;
  wire seg_14_2_neigh_op_tnr_3_56859;
  wire seg_14_2_neigh_op_tnr_7_56863;
  wire seg_14_2_neigh_op_top_3_53029;
  wire seg_14_2_sp12_v_b_12_56584;
  wire seg_14_2_sp4_h_r_10_56870;
  wire seg_14_2_sp4_v_b_14_52911;
  wire seg_14_3_glb_netwk_0_5;
  wire seg_14_3_local_g0_0_56897;
  wire seg_14_3_local_g0_1_56898;
  wire seg_14_3_local_g0_2_56899;
  wire seg_14_3_local_g0_7_56904;
  wire seg_14_3_local_g1_0_56905;
  wire seg_14_3_local_g1_1_56906;
  wire seg_14_3_local_g1_3_56908;
  wire seg_14_3_local_g1_4_56909;
  wire seg_14_3_local_g1_6_56911;
  wire seg_14_3_local_g1_7_56912;
  wire seg_14_3_local_g2_1_56914;
  wire seg_14_3_local_g2_2_56915;
  wire seg_14_3_local_g2_3_56916;
  wire seg_14_3_local_g2_4_56917;
  wire seg_14_3_local_g2_7_56920;
  wire seg_14_3_local_g3_0_56921;
  wire seg_14_3_local_g3_3_56924;
  wire seg_14_3_local_g3_7_56928;
  wire seg_14_3_lutff_0_out_53026;
  wire seg_14_3_lutff_1_out_53027;
  wire seg_14_3_lutff_2_out_53028;
  wire seg_14_3_lutff_3_out_53029;
  wire seg_14_3_lutff_4_out_53030;
  wire seg_14_3_lutff_5_out_53031;
  wire seg_14_3_lutff_6_out_53032;
  wire seg_14_3_lutff_7_out_53033;
  wire seg_14_3_neigh_op_bnr_0_56697;
  wire seg_14_3_neigh_op_bnr_1_56698;
  wire seg_14_3_neigh_op_lft_7_49202;
  wire seg_14_3_neigh_op_rgt_2_56858;
  wire seg_14_3_neigh_op_rgt_3_56859;
  wire seg_14_3_neigh_op_rgt_7_56863;
  wire seg_14_3_neigh_op_top_0_53149;
  wire seg_14_3_neigh_op_top_1_53150;
  wire seg_14_3_neigh_op_top_4_53153;
  wire seg_14_3_neigh_op_top_7_53156;
  wire seg_14_3_sp12_v_b_11_56584;
  wire seg_14_3_sp4_r_v_b_12_56751;
  wire seg_14_3_sp4_v_b_14_52923;
  wire seg_14_3_sp4_v_b_19_52929;
  wire seg_14_3_sp4_v_t_42_53302;
  wire seg_14_4_glb_netwk_0_5;
  wire seg_14_4_local_g0_3_57023;
  wire seg_14_4_local_g0_7_57027;
  wire seg_14_4_local_g1_0_57028;
  wire seg_14_4_local_g1_2_57030;
  wire seg_14_4_local_g1_6_57034;
  wire seg_14_4_local_g2_2_57038;
  wire seg_14_4_local_g2_5_57041;
  wire seg_14_4_local_g3_0_57044;
  wire seg_14_4_local_g3_2_57046;
  wire seg_14_4_local_g3_5_57049;
  wire seg_14_4_local_g3_7_57051;
  wire seg_14_4_lutff_0_out_53149;
  wire seg_14_4_lutff_1_out_53150;
  wire seg_14_4_lutff_2_out_53151;
  wire seg_14_4_lutff_4_out_53153;
  wire seg_14_4_lutff_5_out_53154;
  wire seg_14_4_lutff_7_out_53156;
  wire seg_14_4_neigh_op_bot_0_53026;
  wire seg_14_4_neigh_op_bot_6_53032;
  wire seg_14_4_neigh_op_lft_2_49320;
  wire seg_14_4_neigh_op_lft_3_49321;
  wire seg_14_4_sp4_h_l_36_41792;
  wire seg_14_4_sp4_h_l_41_41797;
  wire seg_14_4_sp4_h_r_29_49460;
  wire seg_14_4_sp4_v_b_42_53302;
  wire seg_14_4_sp4_v_t_38_53421;
  wire seg_14_7_glb_netwk_0_5;
  wire seg_14_7_local_g0_2_57391;
  wire seg_14_7_local_g1_6_57403;
  wire seg_14_7_local_g2_5_57410;
  wire seg_14_7_local_g2_7_57412;
  wire seg_14_7_local_g3_1_57414;
  wire seg_14_7_local_g3_2_57415;
  wire seg_14_7_local_g3_5_57418;
  wire seg_14_7_lutff_1_out_53519;
  wire seg_14_7_lutff_6_out_53524;
  wire seg_14_7_lutff_7_out_53525;
  wire seg_14_7_sp4_h_l_47_42162;
  wire seg_14_7_sp4_h_r_10_57485;
  wire seg_14_7_sp4_h_r_29_49829;
  wire seg_14_7_sp4_h_r_5_57490;
  wire seg_14_7_sp4_h_r_6_57491;
  wire seg_14_7_sp4_r_v_b_18_57255;
  wire seg_14_7_sp4_r_v_b_45_57504;
  wire seg_14_7_sp4_v_b_28_53547;
  wire seg_14_7_sp4_v_t_41_53793;
  wire seg_14_8_glb_netwk_0_5;
  wire seg_14_8_local_g0_3_57515;
  wire seg_14_8_local_g0_6_57518;
  wire seg_14_8_local_g1_3_57523;
  wire seg_14_8_local_g1_6_57526;
  wire seg_14_8_local_g1_7_57527;
  wire seg_14_8_local_g2_0_57528;
  wire seg_14_8_local_g2_1_57529;
  wire seg_14_8_local_g2_7_57535;
  wire seg_14_8_local_g3_0_57536;
  wire seg_14_8_local_g3_3_57539;
  wire seg_14_8_local_g3_5_57541;
  wire seg_14_8_local_g3_7_57543;
  wire seg_14_8_lutff_6_out_53647;
  wire seg_14_8_lutff_7_out_53648;
  wire seg_14_8_neigh_op_bot_6_53524;
  wire seg_14_8_neigh_op_lft_3_49813;
  wire seg_14_8_neigh_op_tnl_0_49933;
  wire seg_14_8_neigh_op_tnl_5_49938;
  wire seg_14_8_neigh_op_top_3_53767;
  wire seg_14_8_neigh_op_top_6_53770;
  wire seg_14_8_sp4_h_l_38_42288;
  wire seg_14_8_sp4_h_r_25_49946;
  wire seg_14_8_sp4_h_r_8_57616;
  wire seg_14_8_sp4_r_v_b_11_57259;
  wire seg_14_8_sp4_r_v_b_25_57495;
  wire seg_14_8_sp4_r_v_b_32_57504;
  wire seg_14_8_sp4_v_b_1_53419;
  wire seg_14_8_sp4_v_b_31_53671;
  wire seg_14_8_sp4_v_b_43_53795;
  wire seg_14_9_local_g0_0_57635;
  wire seg_14_9_local_g0_1_57636;
  wire seg_14_9_local_g0_5_57640;
  wire seg_14_9_local_g0_6_57641;
  wire seg_14_9_local_g0_7_57642;
  wire seg_14_9_local_g1_0_57643;
  wire seg_14_9_local_g1_4_57647;
  wire seg_14_9_local_g1_6_57649;
  wire seg_14_9_local_g2_1_57652;
  wire seg_14_9_local_g3_1_57660;
  wire seg_14_9_lutff_2_out_53766;
  wire seg_14_9_lutff_3_out_53767;
  wire seg_14_9_lutff_4_out_53768;
  wire seg_14_9_lutff_5_out_53769;
  wire seg_14_9_lutff_6_out_53770;
  wire seg_14_9_lutff_7_out_53771;
  wire seg_14_9_neigh_op_bnr_0_57471;
  wire seg_14_9_neigh_op_bot_6_53647;
  wire seg_14_9_neigh_op_bot_7_53648;
  wire seg_14_9_neigh_op_lft_0_49933;
  wire seg_14_9_neigh_op_lft_1_49934;
  wire seg_14_9_neigh_op_lft_5_49938;
  wire seg_14_9_neigh_op_lft_6_49939;
  wire seg_14_9_sp4_v_b_41_53916;
  wire seg_14_9_sp4_v_b_4_53547;
  wire seg_15_0_span4_vert_19_56732;
  wire seg_15_10_glb_netwk_0_5;
  wire seg_15_10_local_g0_0_61588;
  wire seg_15_10_local_g0_3_61591;
  wire seg_15_10_local_g0_4_61592;
  wire seg_15_10_local_g0_6_61594;
  wire seg_15_10_local_g1_0_61596;
  wire seg_15_10_local_g1_2_61598;
  wire seg_15_10_local_g1_3_61599;
  wire seg_15_10_local_g1_4_61600;
  wire seg_15_10_local_g1_5_61601;
  wire seg_15_10_local_g1_6_61602;
  wire seg_15_10_local_g2_5_61609;
  wire seg_15_10_local_g2_6_61610;
  wire seg_15_10_local_g3_1_61613;
  wire seg_15_10_local_g3_4_61616;
  wire seg_15_10_local_g3_5_61617;
  wire seg_15_10_lutff_4_out_57721;
  wire seg_15_10_neigh_op_bnr_6_61430;
  wire seg_15_10_neigh_op_bot_0_57594;
  wire seg_15_10_neigh_op_bot_5_57599;
  wire seg_15_10_neigh_op_rgt_5_61552;
  wire seg_15_10_sp12_v_b_12_60943;
  wire seg_15_10_sp12_v_b_20_61435;
  wire seg_15_10_sp4_h_l_45_46370;
  wire seg_15_10_sp4_h_r_0_61682;
  wire seg_15_10_sp4_h_r_10_61684;
  wire seg_15_10_sp4_h_r_19_57860;
  wire seg_15_10_sp4_h_r_20_57863;
  wire seg_15_10_sp4_h_r_24_54022;
  wire seg_15_10_sp4_h_r_29_54029;
  wire seg_15_10_sp4_h_r_3_61687;
  wire seg_15_10_sp4_h_r_4_61688;
  wire seg_15_10_sp4_h_r_6_61690;
  wire seg_15_10_sp4_h_r_8_61692;
  wire seg_15_10_sp4_r_v_b_17_61453;
  wire seg_15_10_sp4_r_v_b_41_61699;
  wire seg_15_10_sp4_r_v_b_9_61333;
  wire seg_15_10_sp4_v_b_19_57625;
  wire seg_15_10_sp4_v_b_1_57495;
  wire seg_15_10_sp4_v_b_24_57742;
  wire seg_15_10_sp4_v_b_38_57866;
  wire seg_15_10_sp4_v_b_40_57868;
  wire seg_15_10_sp4_v_b_42_57870;
  wire seg_15_11_glb_netwk_0_5;
  wire seg_15_11_local_g0_4_61715;
  wire seg_15_11_local_g0_5_61716;
  wire seg_15_11_local_g0_6_61717;
  wire seg_15_11_local_g1_0_61719;
  wire seg_15_11_local_g1_5_61724;
  wire seg_15_11_local_g1_7_61726;
  wire seg_15_11_local_g2_1_61728;
  wire seg_15_11_local_g2_2_61729;
  wire seg_15_11_local_g2_3_61730;
  wire seg_15_11_local_g2_4_61731;
  wire seg_15_11_local_g3_0_61735;
  wire seg_15_11_local_g3_1_61736;
  wire seg_15_11_local_g3_2_61737;
  wire seg_15_11_local_g3_3_61738;
  wire seg_15_11_local_g3_4_61739;
  wire seg_15_11_local_g3_5_61740;
  wire seg_15_11_local_g3_6_61741;
  wire seg_15_11_lutff_1_out_57841;
  wire seg_15_11_lutff_2_out_57842;
  wire seg_15_11_lutff_4_out_57844;
  wire seg_15_11_lutff_6_out_57846;
  wire seg_15_11_lutff_7_out_57847;
  wire seg_15_11_neigh_op_bnr_5_61552;
  wire seg_15_11_neigh_op_lft_0_54010;
  wire seg_15_11_neigh_op_lft_5_54015;
  wire seg_15_11_neigh_op_lft_6_54016;
  wire seg_15_11_neigh_op_rgt_0_61670;
  wire seg_15_11_neigh_op_rgt_1_61671;
  wire seg_15_11_neigh_op_rgt_4_61674;
  wire seg_15_11_sp12_v_b_10_60942;
  wire seg_15_11_sp4_h_r_22_57978;
  wire seg_15_11_sp4_h_r_37_50314;
  wire seg_15_11_sp4_r_v_b_20_61579;
  wire seg_15_11_sp4_r_v_b_22_61581;
  wire seg_15_11_sp4_r_v_b_27_61696;
  wire seg_15_11_sp4_v_b_15_57744;
  wire seg_15_11_sp4_v_b_20_57749;
  wire seg_15_11_sp4_v_b_33_57872;
  wire seg_15_11_sp4_v_b_34_57875;
  wire seg_15_11_sp4_v_b_35_57874;
  wire seg_15_11_sp4_v_b_43_57994;
  wire seg_15_12_glb_netwk_0_5;
  wire seg_15_12_local_g0_3_61837;
  wire seg_15_12_local_g0_4_61838;
  wire seg_15_12_local_g0_7_61841;
  wire seg_15_12_local_g1_0_61842;
  wire seg_15_12_local_g1_3_61845;
  wire seg_15_12_local_g2_0_61850;
  wire seg_15_12_local_g2_1_61851;
  wire seg_15_12_local_g2_2_61852;
  wire seg_15_12_local_g2_4_61854;
  wire seg_15_12_local_g2_5_61855;
  wire seg_15_12_local_g2_6_61856;
  wire seg_15_12_local_g2_7_61857;
  wire seg_15_12_local_g3_2_61860;
  wire seg_15_12_local_g3_3_61861;
  wire seg_15_12_local_g3_4_61862;
  wire seg_15_12_local_g3_5_61863;
  wire seg_15_12_local_g3_6_61864;
  wire seg_15_12_lutff_0_out_57963;
  wire seg_15_12_lutff_1_out_57964;
  wire seg_15_12_lutff_2_out_57965;
  wire seg_15_12_lutff_3_out_57966;
  wire seg_15_12_lutff_4_out_57967;
  wire seg_15_12_lutff_5_out_57968;
  wire seg_15_12_lutff_6_out_57969;
  wire seg_15_12_lutff_7_out_57970;
  wire seg_15_12_neigh_op_top_3_58089;
  wire seg_15_12_neigh_op_top_4_58090;
  wire seg_15_12_sp4_h_l_37_46606;
  wire seg_15_12_sp4_h_l_38_46611;
  wire seg_15_12_sp4_h_l_41_46612;
  wire seg_15_12_sp4_h_l_45_46616;
  wire seg_15_12_sp4_r_v_b_0_61572;
  wire seg_15_12_sp4_r_v_b_31_61823;
  wire seg_15_12_sp4_v_b_0_57742;
  wire seg_15_12_sp4_v_b_11_57751;
  wire seg_15_12_sp4_v_b_25_57987;
  wire seg_15_12_sp4_v_b_27_57989;
  wire seg_15_12_sp4_v_b_28_57992;
  wire seg_15_12_sp4_v_b_29_57991;
  wire seg_15_12_sp4_v_b_34_57998;
  wire seg_15_12_sp4_v_b_36_58110;
  wire seg_15_12_sp4_v_b_38_58112;
  wire seg_15_12_sp4_v_b_40_58114;
  wire seg_15_12_sp4_v_b_42_58116;
  wire seg_15_12_sp4_v_b_45_58119;
  wire seg_15_12_sp4_v_b_46_58120;
  wire seg_15_12_sp4_v_b_47_58121;
  wire seg_15_12_sp4_v_t_46_58243;
  wire seg_15_12_sp4_v_t_47_58244;
  wire seg_15_13_local_g0_0_61957;
  wire seg_15_13_local_g0_4_61961;
  wire seg_15_13_local_g0_5_61962;
  wire seg_15_13_local_g0_6_61963;
  wire seg_15_13_local_g1_0_61965;
  wire seg_15_13_local_g1_1_61966;
  wire seg_15_13_local_g1_2_61967;
  wire seg_15_13_local_g1_3_61968;
  wire seg_15_13_local_g1_4_61969;
  wire seg_15_13_local_g1_5_61970;
  wire seg_15_13_local_g1_7_61972;
  wire seg_15_13_local_g2_0_61973;
  wire seg_15_13_local_g2_1_61974;
  wire seg_15_13_local_g2_3_61976;
  wire seg_15_13_local_g2_4_61977;
  wire seg_15_13_local_g2_5_61978;
  wire seg_15_13_local_g3_2_61983;
  wire seg_15_13_local_g3_3_61984;
  wire seg_15_13_local_g3_4_61985;
  wire seg_15_13_local_g3_5_61986;
  wire seg_15_13_lutff_3_out_58089;
  wire seg_15_13_lutff_4_out_58090;
  wire seg_15_13_lutff_7_out_58093;
  wire seg_15_13_neigh_op_bot_0_57963;
  wire seg_15_13_neigh_op_bot_2_57965;
  wire seg_15_13_neigh_op_bot_4_57967;
  wire seg_15_13_neigh_op_bot_5_57968;
  wire seg_15_13_neigh_op_tnl_1_54380;
  wire seg_15_13_neigh_op_top_0_58209;
  wire seg_15_13_neigh_op_top_5_58214;
  wire seg_15_13_sp4_h_l_38_46734;
  wire seg_15_13_sp4_h_l_43_46737;
  wire seg_15_13_sp4_h_l_44_46740;
  wire seg_15_13_sp4_h_l_46_46732;
  wire seg_15_13_sp4_h_l_47_46731;
  wire seg_15_13_sp4_h_r_0_62051;
  wire seg_15_13_sp4_h_r_10_62053;
  wire seg_15_13_sp4_h_r_12_58222;
  wire seg_15_13_sp4_h_r_17_58227;
  wire seg_15_13_sp4_h_r_18_58230;
  wire seg_15_13_sp4_h_r_27_54396;
  wire seg_15_13_sp4_h_r_28_54397;
  wire seg_15_13_sp4_h_r_32_54401;
  wire seg_15_13_sp4_h_r_4_62057;
  wire seg_15_13_sp4_r_v_b_13_61818;
  wire seg_15_13_sp4_r_v_b_19_61824;
  wire seg_15_13_sp4_r_v_b_3_61696;
  wire seg_15_13_sp4_r_v_b_4_61699;
  wire seg_15_13_sp4_v_b_26_58113;
  wire seg_15_13_sp4_v_b_2_57867;
  wire seg_15_13_sp4_v_b_36_58233;
  wire seg_15_13_sp4_v_b_37_58234;
  wire seg_15_13_sp4_v_b_43_58240;
  wire seg_15_13_sp4_v_b_45_58242;
  wire seg_15_13_sp4_v_b_6_57871;
  wire seg_15_13_sp4_v_t_37_58357;
  wire seg_15_13_sp4_v_t_38_58358;
  wire seg_15_14_glb_netwk_0_5;
  wire seg_15_14_glb_netwk_3_8;
  wire seg_15_14_local_g0_1_62081;
  wire seg_15_14_local_g0_2_62082;
  wire seg_15_14_local_g0_3_62083;
  wire seg_15_14_local_g0_6_62086;
  wire seg_15_14_local_g1_1_62089;
  wire seg_15_14_local_g1_2_62090;
  wire seg_15_14_local_g1_4_62092;
  wire seg_15_14_local_g1_6_62094;
  wire seg_15_14_local_g1_7_62095;
  wire seg_15_14_local_g2_0_62096;
  wire seg_15_14_local_g2_2_62098;
  wire seg_15_14_local_g2_4_62100;
  wire seg_15_14_local_g2_5_62101;
  wire seg_15_14_local_g3_1_62105;
  wire seg_15_14_local_g3_7_62111;
  wire seg_15_14_lutff_0_out_58209;
  wire seg_15_14_lutff_5_out_58214;
  wire seg_15_14_neigh_op_bnl_2_54258;
  wire seg_15_14_neigh_op_lft_6_54385;
  wire seg_15_14_neigh_op_top_1_58333;
  wire seg_15_14_neigh_op_top_7_58339;
  wire seg_15_14_sp12_v_b_4_60943;
  wire seg_15_14_sp4_h_l_36_46853;
  wire seg_15_14_sp4_h_l_37_46852;
  wire seg_15_14_sp4_h_l_38_46857;
  wire seg_15_14_sp4_h_l_44_46863;
  wire seg_15_14_sp4_h_l_45_46862;
  wire seg_15_14_sp4_h_l_46_46855;
  wire seg_15_14_sp4_h_l_47_46854;
  wire seg_15_14_sp4_h_r_11_62177;
  wire seg_15_14_sp4_h_r_14_58349;
  wire seg_15_14_sp4_h_r_2_62178;
  wire seg_15_14_sp4_h_r_41_50689;
  wire seg_15_14_sp4_h_r_4_62180;
  wire seg_15_14_sp4_h_r_6_62182;
  wire seg_15_14_sp4_h_r_8_62184;
  wire seg_15_14_sp4_r_v_b_15_61943;
  wire seg_15_14_sp4_r_v_b_19_61947;
  wire seg_15_14_sp4_r_v_b_33_62071;
  wire seg_15_14_sp4_r_v_b_7_61823;
  wire seg_15_14_sp4_v_b_0_57988;
  wire seg_15_14_sp4_v_b_12_58110;
  wire seg_15_14_sp4_v_b_1_57987;
  wire seg_15_14_sp4_v_b_2_57990;
  wire seg_15_14_sp4_v_b_47_58367;
  wire seg_15_14_sp4_v_b_4_57992;
  wire seg_15_14_sp4_v_b_7_57993;
  wire seg_15_14_sp4_v_b_8_57996;
  wire seg_15_14_sp4_v_b_9_57995;
  wire seg_15_14_sp4_v_t_46_58489;
  wire seg_15_15_glb_netwk_0_5;
  wire seg_15_15_glb_netwk_3_8;
  wire seg_15_15_local_g0_1_62204;
  wire seg_15_15_local_g0_3_62206;
  wire seg_15_15_local_g0_5_62208;
  wire seg_15_15_local_g0_6_62209;
  wire seg_15_15_local_g0_7_62210;
  wire seg_15_15_local_g1_6_62217;
  wire seg_15_15_local_g1_7_62218;
  wire seg_15_15_local_g2_1_62220;
  wire seg_15_15_local_g2_2_62221;
  wire seg_15_15_local_g2_5_62224;
  wire seg_15_15_local_g3_0_62227;
  wire seg_15_15_local_g3_2_62229;
  wire seg_15_15_local_g3_3_62230;
  wire seg_15_15_local_g3_5_62232;
  wire seg_15_15_lutff_0_out_58332;
  wire seg_15_15_lutff_1_out_58333;
  wire seg_15_15_lutff_5_out_58337;
  wire seg_15_15_lutff_7_out_58339;
  wire seg_15_15_neigh_op_tnl_5_54630;
  wire seg_15_15_sp4_h_l_38_46980;
  wire seg_15_15_sp4_h_l_39_46979;
  wire seg_15_15_sp4_h_l_40_46982;
  wire seg_15_15_sp4_h_l_42_46984;
  wire seg_15_15_sp4_h_l_43_46983;
  wire seg_15_15_sp4_h_l_46_46978;
  wire seg_15_15_sp4_h_r_11_62300;
  wire seg_15_15_sp4_h_r_13_58467;
  wire seg_15_15_sp4_h_r_26_54641;
  wire seg_15_15_sp4_h_r_41_50812;
  wire seg_15_15_sp4_h_r_4_62303;
  wire seg_15_15_sp4_h_r_6_62305;
  wire seg_15_15_sp4_h_r_7_62306;
  wire seg_15_15_sp4_h_r_8_62307;
  wire seg_15_15_sp4_r_v_b_13_62064;
  wire seg_15_15_sp4_r_v_b_31_62192;
  wire seg_15_15_sp4_v_b_14_58235;
  wire seg_15_15_sp4_v_b_22_58243;
  wire seg_15_15_sp4_v_b_26_58359;
  wire seg_15_15_sp4_v_b_35_58366;
  wire seg_15_15_sp4_v_t_43_58609;
  wire seg_15_16_glb_netwk_0_5;
  wire seg_15_16_local_g0_1_62327;
  wire seg_15_16_local_g0_5_62331;
  wire seg_15_16_local_g1_0_62334;
  wire seg_15_16_local_g1_3_62337;
  wire seg_15_16_local_g1_5_62339;
  wire seg_15_16_local_g1_6_62340;
  wire seg_15_16_local_g2_2_62344;
  wire seg_15_16_local_g2_4_62346;
  wire seg_15_16_local_g2_6_62348;
  wire seg_15_16_local_g3_0_62350;
  wire seg_15_16_local_g3_3_62353;
  wire seg_15_16_local_g3_4_62354;
  wire seg_15_16_local_g3_6_62356;
  wire seg_15_16_lutff_6_out_58461;
  wire seg_15_16_neigh_op_rgt_2_62287;
  wire seg_15_16_sp4_h_l_39_47102;
  wire seg_15_16_sp4_h_r_17_58596;
  wire seg_15_16_sp4_h_r_26_54764;
  wire seg_15_16_sp4_h_r_5_62427;
  wire seg_15_16_sp4_h_r_6_62428;
  wire seg_15_16_sp4_r_v_b_20_62194;
  wire seg_15_16_sp4_r_v_b_22_62196;
  wire seg_15_16_sp4_r_v_b_5_62067;
  wire seg_15_16_sp4_r_v_b_9_62071;
  wire seg_15_16_sp4_v_b_0_58234;
  wire seg_15_16_sp4_v_b_14_58358;
  wire seg_15_16_sp4_v_b_16_58360;
  wire seg_15_16_sp4_v_b_19_58363;
  wire seg_15_16_sp4_v_b_28_58484;
  wire seg_15_16_sp4_v_b_2_58236;
  wire seg_15_16_sp4_v_b_32_58488;
  wire seg_15_16_sp4_v_b_3_58235;
  wire seg_15_16_sp4_v_b_43_58609;
  wire seg_15_16_sp4_v_b_5_58237;
  wire seg_15_16_sp4_v_b_6_58240;
  wire seg_15_16_sp4_v_b_9_58241;
  wire seg_15_16_sp4_v_t_37_58726;
  wire seg_15_16_sp4_v_t_38_58727;
  wire seg_15_16_sp4_v_t_46_58735;
  wire seg_15_17_glb_netwk_0_5;
  wire seg_15_17_local_g0_7_62456;
  wire seg_15_17_local_g1_0_62457;
  wire seg_15_17_local_g1_1_62458;
  wire seg_15_17_local_g1_3_62460;
  wire seg_15_17_local_g2_2_62467;
  wire seg_15_17_local_g2_4_62469;
  wire seg_15_17_local_g2_5_62470;
  wire seg_15_17_local_g2_6_62471;
  wire seg_15_17_local_g2_7_62472;
  wire seg_15_17_local_g3_5_62478;
  wire seg_15_17_local_g3_6_62479;
  wire seg_15_17_lutff_0_out_58578;
  wire seg_15_17_lutff_2_out_58580;
  wire seg_15_17_lutff_7_out_58585;
  wire seg_15_17_sp4_h_l_46_47224;
  wire seg_15_17_sp4_h_r_19_58721;
  wire seg_15_17_sp4_h_r_28_54889;
  wire seg_15_17_sp4_h_r_29_54890;
  wire seg_15_17_sp4_h_r_7_62552;
  wire seg_15_17_sp4_r_v_b_12_62309;
  wire seg_15_17_sp4_r_v_b_22_62319;
  wire seg_15_17_sp4_v_b_10_58367;
  wire seg_15_17_sp4_v_b_17_58484;
  wire seg_15_17_sp4_v_b_22_58489;
  wire seg_15_17_sp4_v_b_2_58359;
  wire seg_15_17_sp4_v_b_30_58609;
  wire seg_15_17_sp4_v_b_37_58726;
  wire seg_15_17_sp4_v_t_38_58850;
  wire seg_15_17_sp4_v_t_40_58852;
  wire seg_15_17_sp4_v_t_41_58853;
  wire seg_15_17_sp4_v_t_44_58856;
  wire seg_15_18_glb_netwk_0_5;
  wire seg_15_18_glb_netwk_3_8;
  wire seg_15_18_local_g0_0_62572;
  wire seg_15_18_local_g0_1_62573;
  wire seg_15_18_local_g0_2_62574;
  wire seg_15_18_local_g0_6_62578;
  wire seg_15_18_local_g0_7_62579;
  wire seg_15_18_local_g1_2_62582;
  wire seg_15_18_local_g1_4_62584;
  wire seg_15_18_local_g2_0_62588;
  wire seg_15_18_local_g2_1_62589;
  wire seg_15_18_local_g2_4_62592;
  wire seg_15_18_local_g2_5_62593;
  wire seg_15_18_local_g3_1_62597;
  wire seg_15_18_local_g3_3_62599;
  wire seg_15_18_local_g3_4_62600;
  wire seg_15_18_lutff_1_out_58702;
  wire seg_15_18_lutff_2_out_58703;
  wire seg_15_18_lutff_4_out_58705;
  wire seg_15_18_lutff_7_out_58708;
  wire seg_15_18_neigh_op_tnl_1_54995;
  wire seg_15_18_neigh_op_top_0_58824;
  wire seg_15_18_neigh_op_top_6_58830;
  wire seg_15_18_sp12_h_r_0_62662;
  wire seg_15_18_sp4_h_l_39_47348;
  wire seg_15_18_sp4_h_l_40_47351;
  wire seg_15_18_sp4_h_r_0_62666;
  wire seg_15_18_sp4_h_r_12_58837;
  wire seg_15_18_sp4_h_r_25_55007;
  wire seg_15_18_sp4_h_r_2_62670;
  wire seg_15_18_sp4_h_r_35_55009;
  wire seg_15_18_sp4_r_v_b_12_62432;
  wire seg_15_18_sp4_r_v_b_13_62433;
  wire seg_15_18_sp4_v_b_10_58490;
  wire seg_15_18_sp4_v_b_24_58726;
  wire seg_15_18_sp4_v_b_4_58484;
  wire seg_15_18_sp4_v_t_36_58971;
  wire seg_15_18_sp4_v_t_38_58973;
  wire seg_15_18_sp4_v_t_45_58980;
  wire seg_15_19_glb_netwk_0_5;
  wire seg_15_19_local_g0_7_62702;
  wire seg_15_19_local_g1_0_62703;
  wire seg_15_19_local_g1_3_62706;
  wire seg_15_19_local_g2_4_62715;
  wire seg_15_19_local_g3_1_62720;
  wire seg_15_19_local_g3_3_62722;
  wire seg_15_19_local_g3_4_62723;
  wire seg_15_19_local_g3_5_62724;
  wire seg_15_19_lutff_0_out_58824;
  wire seg_15_19_lutff_3_out_58827;
  wire seg_15_19_lutff_5_out_58829;
  wire seg_15_19_lutff_6_out_58830;
  wire seg_15_19_neigh_op_top_0_58947;
  wire seg_15_19_sp4_h_l_45_47477;
  wire seg_15_19_sp4_h_r_22_58962;
  wire seg_15_19_sp4_h_r_23_58961;
  wire seg_15_19_sp4_h_r_28_55135;
  wire seg_15_19_sp4_h_r_38_51303;
  wire seg_15_19_sp4_h_r_6_62797;
  wire seg_15_19_sp4_r_v_b_20_62563;
  wire seg_15_19_sp4_r_v_b_23_62566;
  wire seg_15_19_sp4_r_v_b_27_62680;
  wire seg_15_19_sp4_r_v_b_7_62438;
  wire seg_15_19_sp4_v_b_22_58735;
  wire seg_15_19_sp4_v_b_33_58856;
  wire seg_15_19_sp4_v_b_6_58609;
  wire seg_15_20_glb_netwk_0_5;
  wire seg_15_20_local_g0_0_62818;
  wire seg_15_20_local_g0_3_62821;
  wire seg_15_20_local_g1_2_62828;
  wire seg_15_20_local_g1_3_62829;
  wire seg_15_20_local_g1_7_62833;
  wire seg_15_20_local_g2_0_62834;
  wire seg_15_20_local_g2_4_62838;
  wire seg_15_20_local_g3_2_62844;
  wire seg_15_20_local_g3_7_62849;
  wire seg_15_20_lutff_0_out_58947;
  wire seg_15_20_lutff_2_out_58949;
  wire seg_15_20_neigh_op_bot_3_58827;
  wire seg_15_20_sp12_v_b_0_61435;
  wire seg_15_20_sp4_h_l_36_47591;
  wire seg_15_20_sp4_h_l_47_47592;
  wire seg_15_20_sp4_h_r_30_55260;
  wire seg_15_20_sp4_h_r_44_51432;
  wire seg_15_20_sp4_h_r_8_62922;
  wire seg_15_20_sp4_r_v_b_18_62684;
  wire seg_15_20_sp4_r_v_b_1_62555;
  wire seg_15_20_sp4_r_v_b_36_62924;
  wire seg_15_20_sp4_r_v_b_3_62557;
  wire seg_15_20_sp4_r_v_b_7_62561;
  wire seg_15_20_sp4_v_b_0_58726;
  wire seg_15_20_sp4_v_b_14_58850;
  wire seg_15_20_sp4_v_b_16_58852;
  wire seg_15_20_sp4_v_b_40_59098;
  wire seg_15_20_sp4_v_b_47_59105;
  wire seg_15_20_sp4_v_t_37_59218;
  wire seg_15_20_sp4_v_t_38_59219;
  wire seg_15_21_local_g1_7_62956;
  wire seg_15_21_local_g3_2_62967;
  wire seg_15_21_sp4_h_l_38_47718;
  wire seg_15_21_sp4_h_l_44_47724;
  wire seg_15_21_sp4_h_r_12_59206;
  wire seg_15_21_sp4_h_r_28_55381;
  wire seg_15_21_sp4_h_r_3_63040;
  wire seg_15_21_sp4_h_r_44_51555;
  wire seg_15_21_sp4_r_v_b_13_62802;
  wire seg_15_21_sp4_r_v_b_7_62684;
  wire seg_15_21_sp4_v_b_12_58971;
  wire seg_15_21_sp4_v_b_34_59105;
  wire seg_15_22_glb_netwk_0_5;
  wire seg_15_22_local_g0_4_63068;
  wire seg_15_22_local_g1_7_63079;
  wire seg_15_22_local_g3_3_63091;
  wire seg_15_22_lutff_4_out_59197;
  wire seg_15_22_lutff_5_out_59198;
  wire seg_15_22_sp4_h_r_23_59330;
  wire seg_15_22_sp4_r_v_b_19_62931;
  wire seg_15_22_sp4_v_b_24_59218;
  wire seg_15_22_sp4_v_b_8_58980;
  wire seg_15_23_glb_netwk_0_5;
  wire seg_15_23_local_g0_4_63191;
  wire seg_15_23_local_g0_5_63192;
  wire seg_15_23_local_g1_5_63200;
  wire seg_15_23_local_g2_1_63204;
  wire seg_15_23_local_g2_2_63205;
  wire seg_15_23_lutff_1_out_59317;
  wire seg_15_23_neigh_op_bot_5_59198;
  wire seg_15_23_sp4_h_r_12_59452;
  wire seg_15_23_sp4_h_r_13_59451;
  wire seg_15_23_sp4_h_r_42_51799;
  wire seg_15_23_sp4_v_b_10_59105;
  wire seg_15_23_sp4_v_b_14_59219;
  wire seg_15_23_sp4_v_b_34_59351;
  wire seg_15_23_sp4_v_t_39_59589;
  wire seg_15_25_glb_netwk_0_5;
  wire seg_15_25_local_g0_6_63439;
  wire seg_15_25_local_g1_3_63444;
  wire seg_15_25_sp12_h_r_14_36709;
  wire seg_15_25_sp4_r_v_b_11_63180;
  wire seg_15_25_sp4_r_v_b_27_63418;
  wire seg_15_25_sp4_v_b_10_59351;
  wire seg_15_25_sp4_v_b_26_59589;
  wire seg_15_25_sp4_v_b_3_59342;
  wire seg_15_25_sp4_v_t_42_59838;
  wire seg_15_27_local_g0_4_63683;
  wire seg_15_27_local_g3_7_63710;
  wire seg_15_27_neigh_op_top_4_59935;
  wire seg_15_27_sp12_v_b_7_62665;
  wire seg_15_27_sp4_v_b_10_59597;
  wire seg_15_28_local_g0_5_63807;
  wire seg_15_28_local_g2_1_63819;
  wire seg_15_28_local_g2_5_63823;
  wire seg_15_28_local_g2_6_63824;
  wire seg_15_28_local_g3_3_63829;
  wire seg_15_28_local_g3_4_63830;
  wire seg_15_28_local_g3_5_63831;
  wire seg_15_28_lutff_0_out_59931;
  wire seg_15_28_lutff_4_out_59935;
  wire seg_15_28_lutff_5_out_59936;
  wire seg_15_28_neigh_op_rgt_1_63762;
  wire seg_15_28_neigh_op_rgt_3_63764;
  wire seg_15_28_neigh_op_rgt_5_63766;
  wire seg_15_28_neigh_op_rgt_6_63767;
  wire seg_15_28_sp12_v_b_4_62665;
  wire seg_15_28_sp4_h_l_42_48583;
  wire seg_15_28_sp4_h_r_30_56244;
  wire seg_15_28_sp4_h_r_46_52408;
  wire seg_15_28_sp4_v_b_18_59838;
  wire seg_15_28_sp4_v_b_1_59709;
  wire seg_15_29_local_g0_3_63928;
  wire seg_15_29_local_g0_5_63930;
  wire seg_15_29_local_g1_1_63934;
  wire seg_15_29_local_g1_3_63936;
  wire seg_15_29_local_g1_5_63938;
  wire seg_15_29_local_g1_6_63939;
  wire seg_15_29_local_g3_5_63954;
  wire seg_15_29_lutff_5_out_60059;
  wire seg_15_29_neigh_op_bnr_1_63762;
  wire seg_15_29_neigh_op_bnr_3_63764;
  wire seg_15_29_neigh_op_bnr_5_63766;
  wire seg_15_29_neigh_op_bnr_6_63767;
  wire seg_15_29_sp4_r_v_b_31_63914;
  wire seg_15_29_sp4_v_b_11_59842;
  wire seg_15_2_glb_netwk_0_5;
  wire seg_15_2_local_g0_0_60604;
  wire seg_15_2_local_g0_2_60606;
  wire seg_15_2_local_g0_6_60610;
  wire seg_15_2_local_g0_7_60611;
  wire seg_15_2_local_g1_2_60614;
  wire seg_15_2_local_g1_3_60615;
  wire seg_15_2_local_g3_0_60628;
  wire seg_15_2_lutff_0_out_56697;
  wire seg_15_2_lutff_1_out_56698;
  wire seg_15_2_lutff_2_out_56699;
  wire seg_15_2_lutff_6_out_56703;
  wire seg_15_2_neigh_op_top_2_56858;
  wire seg_15_2_neigh_op_top_3_56859;
  wire seg_15_2_neigh_op_top_7_56863;
  wire seg_15_2_sp4_r_v_b_16_60573;
  wire seg_15_2_sp4_v_b_6_56732;
  wire seg_15_30_sp4_h_l_43_48824;
  wire seg_15_31_span4_vert_43_64169;
  wire seg_15_3_glb_netwk_0_5;
  wire seg_15_3_local_g0_2_60729;
  wire seg_15_3_local_g0_5_60732;
  wire seg_15_3_local_g1_0_60735;
  wire seg_15_3_local_g1_1_60736;
  wire seg_15_3_local_g1_3_60738;
  wire seg_15_3_local_g1_4_60739;
  wire seg_15_3_local_g1_5_60740;
  wire seg_15_3_local_g2_4_60747;
  wire seg_15_3_local_g2_6_60749;
  wire seg_15_3_local_g3_2_60753;
  wire seg_15_3_local_g3_3_60754;
  wire seg_15_3_local_g3_7_60758;
  wire seg_15_3_lutff_1_out_56857;
  wire seg_15_3_lutff_2_out_56858;
  wire seg_15_3_lutff_3_out_56859;
  wire seg_15_3_lutff_4_out_56860;
  wire seg_15_3_lutff_6_out_56862;
  wire seg_15_3_lutff_7_out_56863;
  wire seg_15_3_neigh_op_bnr_5_60532;
  wire seg_15_3_neigh_op_bot_0_56697;
  wire seg_15_3_neigh_op_bot_2_56699;
  wire seg_15_3_neigh_op_lft_4_53030;
  wire seg_15_3_neigh_op_lft_5_53031;
  wire seg_15_3_sp4_h_r_35_53164;
  wire seg_15_3_sp4_r_v_b_43_60840;
  wire seg_15_4_sp4_h_l_42_45631;
  wire seg_15_6_glb_netwk_0_5;
  wire seg_15_6_local_g2_7_61119;
  wire seg_15_6_local_g3_3_61123;
  wire seg_15_6_sp4_h_r_36_49700;
  wire seg_15_6_sp4_h_r_43_49707;
  wire seg_15_6_sp4_r_v_b_21_60965;
  wire seg_15_6_sp4_r_v_b_37_61203;
  wire seg_15_6_sp4_v_b_31_57255;
  wire seg_15_8_glb_netwk_0_5;
  wire seg_15_8_local_g1_0_61350;
  wire seg_15_8_local_g1_3_61353;
  wire seg_15_8_lutff_0_out_57471;
  wire seg_15_8_sp4_h_r_32_53786;
  wire seg_15_8_sp4_r_v_b_17_61207;
  wire seg_15_8_sp4_v_b_11_57259;
  wire seg_15_9_glb_netwk_0_5;
  wire seg_15_9_local_g1_0_61473;
  wire seg_15_9_local_g1_3_61476;
  wire seg_15_9_local_g2_2_61483;
  wire seg_15_9_local_g2_4_61485;
  wire seg_15_9_local_g2_5_61486;
  wire seg_15_9_lutff_0_out_57594;
  wire seg_15_9_lutff_5_out_57599;
  wire seg_15_9_neigh_op_rgt_2_61426;
  wire seg_15_9_neigh_op_rgt_5_61429;
  wire seg_15_9_sp12_v_b_14_60942;
  wire seg_15_9_sp12_v_b_23_61435;
  wire seg_15_9_sp4_r_v_b_0_61203;
  wire seg_15_9_sp4_r_v_b_36_61571;
  wire seg_15_9_sp4_v_b_30_57625;
  wire seg_15_9_sp4_v_b_3_57374;
  wire seg_15_9_sp4_v_b_46_57751;
  wire seg_15_9_sp4_v_t_42_57870;
  wire seg_16_10_local_g1_1_65428;
  wire seg_16_10_lutff_5_out_61552;
  wire seg_16_10_neigh_op_bnr_1_65256;
  wire seg_16_10_sp4_v_b_9_61333;
  wire seg_16_11_glb_netwk_0_5;
  wire seg_16_11_glb_netwk_3_8;
  wire seg_16_11_local_g0_5_65547;
  wire seg_16_11_local_g0_6_65548;
  wire seg_16_11_local_g1_2_65552;
  wire seg_16_11_local_g3_0_65566;
  wire seg_16_11_lutff_0_out_61670;
  wire seg_16_11_lutff_1_out_61671;
  wire seg_16_11_lutff_4_out_61674;
  wire seg_16_11_lutff_5_out_61675;
  wire seg_16_11_neigh_op_top_2_61795;
  wire seg_16_11_sp4_r_v_b_16_65406;
  wire seg_16_11_sp4_v_b_22_61581;
  wire seg_16_12_glb_netwk_0_5;
  wire seg_16_12_glb_netwk_3_8;
  wire seg_16_12_local_g0_2_65667;
  wire seg_16_12_local_g1_1_65674;
  wire seg_16_12_local_g1_2_65675;
  wire seg_16_12_local_g1_4_65677;
  wire seg_16_12_local_g1_5_65678;
  wire seg_16_12_local_g1_6_65679;
  wire seg_16_12_local_g1_7_65680;
  wire seg_16_12_local_g2_2_65683;
  wire seg_16_12_local_g2_3_65684;
  wire seg_16_12_local_g2_5_65686;
  wire seg_16_12_local_g2_6_65687;
  wire seg_16_12_local_g2_7_65688;
  wire seg_16_12_local_g3_0_65689;
  wire seg_16_12_local_g3_4_65693;
  wire seg_16_12_local_g3_6_65695;
  wire seg_16_12_lutff_2_out_61795;
  wire seg_16_12_neigh_op_bnl_4_57844;
  wire seg_16_12_neigh_op_bnl_6_57846;
  wire seg_16_12_neigh_op_bot_5_61675;
  wire seg_16_12_neigh_op_top_4_61920;
  wire seg_16_12_sp4_h_l_36_50438;
  wire seg_16_12_sp4_h_l_40_50444;
  wire seg_16_12_sp4_h_l_42_50446;
  wire seg_16_12_sp4_h_l_46_50440;
  wire seg_16_12_sp4_h_r_0_65759;
  wire seg_16_12_sp4_h_r_12_61929;
  wire seg_16_12_sp4_h_r_14_61933;
  wire seg_16_12_sp4_h_r_18_61937;
  wire seg_16_12_sp4_h_r_26_58102;
  wire seg_16_12_sp4_h_r_2_65763;
  wire seg_16_12_sp4_h_r_40_54275;
  wire seg_16_12_sp4_h_r_43_54276;
  wire seg_16_12_sp4_h_r_47_54270;
  wire seg_16_12_sp4_r_v_b_16_65529;
  wire seg_16_12_sp4_r_v_b_35_65658;
  wire seg_16_12_sp4_v_b_15_61697;
  wire seg_16_12_sp4_v_b_17_61699;
  wire seg_16_12_sp4_v_b_32_61826;
  wire seg_16_12_sp4_v_b_38_61942;
  wire seg_16_12_sp4_v_b_42_61946;
  wire seg_16_12_sp4_v_b_45_61949;
  wire seg_16_12_sp4_v_b_5_61575;
  wire seg_16_12_sp4_v_t_37_62064;
  wire seg_16_12_sp4_v_t_39_62066;
  wire seg_16_13_glb_netwk_0_5;
  wire seg_16_13_local_g0_2_65790;
  wire seg_16_13_local_g0_3_65791;
  wire seg_16_13_local_g0_4_65792;
  wire seg_16_13_local_g1_5_65801;
  wire seg_16_13_local_g2_2_65806;
  wire seg_16_13_local_g2_3_65807;
  wire seg_16_13_local_g3_0_65812;
  wire seg_16_13_local_g3_2_65814;
  wire seg_16_13_lutff_0_out_61916;
  wire seg_16_13_lutff_2_out_61918;
  wire seg_16_13_lutff_3_out_61919;
  wire seg_16_13_lutff_4_out_61920;
  wire seg_16_13_neigh_op_bnl_3_57966;
  wire seg_16_13_neigh_op_top_5_62044;
  wire seg_16_13_sp4_h_l_37_50560;
  wire seg_16_13_sp4_h_l_39_50564;
  wire seg_16_13_sp4_h_l_40_50567;
  wire seg_16_13_sp4_h_r_19_62059;
  wire seg_16_13_sp4_h_r_24_58221;
  wire seg_16_13_sp4_h_r_26_58225;
  wire seg_16_13_sp4_h_r_4_65888;
  wire seg_16_13_sp4_v_b_34_61951;
  wire seg_16_13_sp4_v_b_4_61699;
  wire seg_16_13_sp4_v_t_43_62193;
  wire seg_16_14_glb_netwk_0_5;
  wire seg_16_14_glb_netwk_1_6;
  wire seg_16_14_local_g0_6_65917;
  wire seg_16_14_local_g0_7_65918;
  wire seg_16_14_local_g3_0_65935;
  wire seg_16_14_local_g3_2_65937;
  wire seg_16_14_local_g3_7_65942;
  wire seg_16_14_lutff_1_out_62040;
  wire seg_16_14_lutff_5_out_62044;
  wire seg_16_14_lutff_7_out_62046;
  wire seg_16_14_sp4_h_r_14_62179;
  wire seg_16_14_sp4_v_b_0_61818;
  wire seg_16_14_sp4_v_b_14_61942;
  wire seg_16_14_sp4_v_b_23_61951;
  wire seg_16_14_sp4_v_b_26_62066;
  wire seg_16_14_sp4_v_b_40_62190;
  wire seg_16_14_sp4_v_b_6_61824;
  wire seg_16_14_sp4_v_b_8_61826;
  wire seg_16_14_sp4_v_b_9_61825;
  wire seg_16_14_sp4_v_t_47_62320;
  wire seg_16_15_glb_netwk_0_5;
  wire seg_16_15_glb_netwk_3_8;
  wire seg_16_15_local_g0_0_66034;
  wire seg_16_15_local_g0_1_66035;
  wire seg_16_15_local_g0_2_66036;
  wire seg_16_15_local_g0_6_66040;
  wire seg_16_15_local_g0_7_66041;
  wire seg_16_15_local_g1_0_66042;
  wire seg_16_15_local_g1_7_66049;
  wire seg_16_15_local_g2_0_66050;
  wire seg_16_15_local_g2_4_66054;
  wire seg_16_15_local_g2_5_66055;
  wire seg_16_15_local_g2_6_66056;
  wire seg_16_15_local_g2_7_66057;
  wire seg_16_15_local_g3_3_66061;
  wire seg_16_15_local_g3_4_66062;
  wire seg_16_15_local_g3_7_66065;
  wire seg_16_15_lutff_0_out_62162;
  wire seg_16_15_lutff_3_out_62165;
  wire seg_16_15_lutff_7_out_62169;
  wire seg_16_15_neigh_op_bot_1_62040;
  wire seg_16_15_neigh_op_lft_7_58339;
  wire seg_16_15_neigh_op_top_2_62287;
  wire seg_16_15_sp4_h_l_38_50811;
  wire seg_16_15_sp4_h_l_40_50813;
  wire seg_16_15_sp4_h_r_0_66128;
  wire seg_16_15_sp4_h_r_10_66130;
  wire seg_16_15_sp4_h_r_12_62298;
  wire seg_16_15_sp4_h_r_28_58473;
  wire seg_16_15_sp4_h_r_38_54642;
  wire seg_16_15_sp4_h_r_4_66134;
  wire seg_16_15_sp4_r_v_b_13_65895;
  wire seg_16_15_sp4_r_v_b_15_65897;
  wire seg_16_15_sp4_r_v_b_21_65903;
  wire seg_16_15_sp4_r_v_b_24_66018;
  wire seg_16_15_sp4_v_b_14_62065;
  wire seg_16_15_sp4_v_b_26_62189;
  wire seg_16_15_sp4_v_b_28_62191;
  wire seg_16_15_sp4_v_b_2_61943;
  wire seg_16_15_sp4_v_b_31_62192;
  wire seg_16_15_sp4_v_b_6_61947;
  wire seg_16_15_sp4_v_b_7_61946;
  wire seg_16_15_sp4_v_b_8_61949;
  wire seg_16_15_sp4_v_t_42_62438;
  wire seg_16_16_glb_netwk_0_5;
  wire seg_16_16_local_g0_1_66158;
  wire seg_16_16_local_g2_5_66178;
  wire seg_16_16_local_g3_0_66181;
  wire seg_16_16_local_g3_3_66184;
  wire seg_16_16_lutff_1_out_62286;
  wire seg_16_16_lutff_2_out_62287;
  wire seg_16_16_sp12_v_b_1_64773;
  wire seg_16_16_sp4_h_l_41_50935;
  wire seg_16_16_sp4_h_l_44_50940;
  wire seg_16_16_sp4_h_l_47_50931;
  wire seg_16_16_sp4_h_r_2_66255;
  wire seg_16_16_sp4_h_r_3_66256;
  wire seg_16_16_sp4_r_v_b_13_66018;
  wire seg_16_16_sp4_r_v_b_16_66021;
  wire seg_16_16_sp4_r_v_b_19_66024;
  wire seg_16_16_sp4_v_b_1_62063;
  wire seg_16_16_sp4_v_b_27_62311;
  wire seg_16_16_sp4_v_b_2_62066;
  wire seg_16_16_sp4_v_b_34_62320;
  wire seg_16_16_sp4_v_b_7_62069;
  wire seg_16_16_sp4_v_t_36_62555;
  wire seg_16_16_sp4_v_t_47_62566;
  wire seg_16_17_glb_netwk_0_5;
  wire seg_16_17_glb_netwk_5_10;
  wire seg_16_17_local_g0_1_66281;
  wire seg_16_17_lutff_1_out_62409;
  wire seg_16_17_sp4_h_l_37_51052;
  wire seg_16_17_sp4_h_l_40_51059;
  wire seg_16_17_sp4_h_l_44_51063;
  wire seg_16_17_sp4_h_l_46_51055;
  wire seg_16_17_sp4_h_l_47_51054;
  wire seg_16_17_sp4_v_b_17_62314;
  wire seg_16_17_sp4_v_b_2_62189;
  wire seg_16_17_sp4_v_b_7_62192;
  wire seg_16_18_glb_netwk_0_5;
  wire seg_16_18_local_g0_2_66405;
  wire seg_16_18_local_g0_5_66408;
  wire seg_16_18_local_g1_3_66414;
  wire seg_16_18_local_g1_4_66415;
  wire seg_16_18_local_g1_5_66416;
  wire seg_16_18_local_g2_3_66422;
  wire seg_16_18_local_g3_3_66430;
  wire seg_16_18_local_g3_6_66433;
  wire seg_16_18_lutff_2_out_62533;
  wire seg_16_18_lutff_3_out_62534;
  wire seg_16_18_lutff_4_out_62535;
  wire seg_16_18_neigh_op_lft_2_58703;
  wire seg_16_18_neigh_op_tnl_3_58827;
  wire seg_16_18_neigh_op_top_5_62659;
  wire seg_16_18_sp4_h_l_36_51176;
  wire seg_16_18_sp4_h_l_37_51175;
  wire seg_16_18_sp4_h_l_41_51181;
  wire seg_16_18_sp4_h_l_46_51178;
  wire seg_16_18_sp4_h_r_19_62674;
  wire seg_16_18_sp4_h_r_1_66498;
  wire seg_16_18_sp4_h_r_46_55009;
  wire seg_16_18_sp4_h_r_4_66503;
  wire seg_16_18_sp4_v_b_5_62313;
  wire seg_16_18_sp4_v_t_37_62802;
  wire seg_16_19_glb_netwk_0_5;
  wire seg_16_19_glb_netwk_1_6;
  wire seg_16_19_local_g0_1_66527;
  wire seg_16_19_local_g0_2_66528;
  wire seg_16_19_local_g0_5_66531;
  wire seg_16_19_local_g0_7_66533;
  wire seg_16_19_local_g1_3_66537;
  wire seg_16_19_local_g1_4_66538;
  wire seg_16_19_local_g2_1_66543;
  wire seg_16_19_local_g2_4_66546;
  wire seg_16_19_local_g3_3_66553;
  wire seg_16_19_local_g3_4_66554;
  wire seg_16_19_local_g3_7_66557;
  wire seg_16_19_lutff_1_out_62655;
  wire seg_16_19_lutff_3_out_62657;
  wire seg_16_19_lutff_4_out_62658;
  wire seg_16_19_lutff_5_out_62659;
  wire seg_16_19_lutff_6_out_62660;
  wire seg_16_19_lutff_7_out_62661;
  wire seg_16_19_neigh_op_top_2_62779;
  wire seg_16_19_neigh_op_top_7_62784;
  wire seg_16_19_sp4_h_l_36_51299;
  wire seg_16_19_sp4_h_l_37_51298;
  wire seg_16_19_sp4_h_l_41_51304;
  wire seg_16_19_sp4_h_l_42_51307;
  wire seg_16_19_sp4_h_r_17_62795;
  wire seg_16_19_sp4_h_r_33_58970;
  wire seg_16_19_sp4_h_r_43_55137;
  wire seg_16_19_sp4_v_b_20_62563;
  wire seg_16_19_sp4_v_b_21_62564;
  wire seg_16_19_sp4_v_b_28_62683;
  wire seg_16_20_glb_netwk_0_5;
  wire seg_16_20_local_g0_1_66650;
  wire seg_16_20_local_g0_3_66652;
  wire seg_16_20_local_g0_4_66653;
  wire seg_16_20_local_g0_7_66656;
  wire seg_16_20_local_g1_1_66658;
  wire seg_16_20_local_g1_3_66660;
  wire seg_16_20_local_g1_4_66661;
  wire seg_16_20_local_g1_7_66664;
  wire seg_16_20_local_g2_2_66667;
  wire seg_16_20_local_g3_1_66674;
  wire seg_16_20_local_g3_2_66675;
  wire seg_16_20_local_g3_3_66676;
  wire seg_16_20_lutff_1_out_62778;
  wire seg_16_20_lutff_2_out_62779;
  wire seg_16_20_lutff_3_out_62780;
  wire seg_16_20_lutff_4_out_62781;
  wire seg_16_20_lutff_5_out_62782;
  wire seg_16_20_lutff_7_out_62784;
  wire seg_16_20_neigh_op_rgt_2_66610;
  wire seg_16_20_neigh_op_top_7_62907;
  wire seg_16_20_sp4_h_l_44_51432;
  wire seg_16_20_sp4_h_r_19_62920;
  wire seg_16_20_sp4_h_r_20_62923;
  wire seg_16_20_sp4_h_r_26_59086;
  wire seg_16_20_sp4_r_v_b_43_66762;
  wire seg_16_20_sp4_v_b_10_62566;
  wire seg_16_20_sp4_v_b_17_62683;
  wire seg_16_20_sp4_v_b_19_62685;
  wire seg_16_20_sp4_v_b_23_62689;
  wire seg_16_20_sp4_v_b_9_62563;
  wire seg_16_21_glb_netwk_0_5;
  wire seg_16_21_glb_netwk_1_6;
  wire seg_16_21_local_g3_1_66797;
  wire seg_16_21_lutff_7_out_62907;
  wire seg_16_21_sp4_h_l_37_51544;
  wire seg_16_21_sp4_h_l_41_51550;
  wire seg_16_21_sp4_h_l_44_51555;
  wire seg_16_21_sp4_r_v_b_41_66883;
  wire seg_16_21_sp4_v_t_46_63180;
  wire seg_16_22_sp4_v_b_1_62801;
  wire seg_16_23_sp4_h_l_42_51799;
  wire seg_16_23_sp4_v_t_38_63418;
  wire seg_16_26_sp4_v_b_4_63298;
  wire seg_16_28_glb_netwk_0_5;
  wire seg_16_28_local_g0_0_67633;
  wire seg_16_28_local_g0_2_67635;
  wire seg_16_28_local_g0_4_67637;
  wire seg_16_28_local_g1_1_67642;
  wire seg_16_28_local_g1_2_67643;
  wire seg_16_28_local_g1_4_67645;
  wire seg_16_28_local_g1_6_67647;
  wire seg_16_28_local_g2_0_67649;
  wire seg_16_28_local_g2_1_67650;
  wire seg_16_28_local_g2_5_67654;
  wire seg_16_28_local_g2_7_67656;
  wire seg_16_28_local_g3_0_67657;
  wire seg_16_28_local_g3_3_67660;
  wire seg_16_28_lutff_1_out_63762;
  wire seg_16_28_lutff_2_out_63763;
  wire seg_16_28_lutff_3_out_63764;
  wire seg_16_28_lutff_5_out_63766;
  wire seg_16_28_lutff_6_out_63767;
  wire seg_16_28_lutff_7_out_63768;
  wire seg_16_28_neigh_op_top_0_63884;
  wire seg_16_28_neigh_op_top_4_63888;
  wire seg_16_28_sp12_v_b_1_66249;
  wire seg_16_28_sp4_h_r_12_63897;
  wire seg_16_28_sp4_h_r_24_60066;
  wire seg_16_28_sp4_h_r_2_67731;
  wire seg_16_28_sp4_r_v_b_16_67497;
  wire seg_16_28_sp4_v_b_8_63548;
  wire seg_16_29_glb_netwk_0_5;
  wire seg_16_29_local_g0_1_67757;
  wire seg_16_29_local_g0_2_67758;
  wire seg_16_29_local_g0_3_67759;
  wire seg_16_29_local_g0_5_67761;
  wire seg_16_29_local_g1_1_67765;
  wire seg_16_29_local_g1_3_67767;
  wire seg_16_29_local_g1_6_67770;
  wire seg_16_29_local_g2_0_67772;
  wire seg_16_29_local_g2_2_67774;
  wire seg_16_29_local_g2_6_67778;
  wire seg_16_29_lutff_0_out_63884;
  wire seg_16_29_lutff_2_out_63886;
  wire seg_16_29_lutff_4_out_63888;
  wire seg_16_29_lutff_6_out_63890;
  wire seg_16_29_neigh_op_bot_1_63762;
  wire seg_16_29_neigh_op_bot_3_63764;
  wire seg_16_29_neigh_op_bot_5_63766;
  wire seg_16_29_neigh_op_bot_6_63767;
  wire seg_16_29_sp4_r_v_b_32_67748;
  wire seg_16_29_sp4_v_b_18_63791;
  wire seg_16_2_glb_netwk_0_5;
  wire seg_16_2_local_g0_1_64436;
  wire seg_16_2_local_g1_0_64443;
  wire seg_16_2_local_g1_1_64444;
  wire seg_16_2_local_g1_6_64449;
  wire seg_16_2_local_g2_4_64455;
  wire seg_16_2_local_g2_7_64458;
  wire seg_16_2_local_g3_2_64461;
  wire seg_16_2_local_g3_3_64462;
  wire seg_16_2_local_g3_7_64466;
  wire seg_16_2_lutff_1_out_60528;
  wire seg_16_2_lutff_2_out_60529;
  wire seg_16_2_lutff_5_out_60532;
  wire seg_16_2_neigh_op_lft_0_56697;
  wire seg_16_2_neigh_op_lft_1_56698;
  wire seg_16_2_neigh_op_lft_6_56703;
  wire seg_16_2_neigh_op_tnl_7_56863;
  wire seg_16_2_sp4_h_r_6_64537;
  wire seg_16_2_sp4_r_v_b_12_64400;
  wire seg_16_2_sp4_r_v_b_19_64406;
  wire seg_16_31_span4_vert_7_63914;
  wire seg_16_3_sp4_h_l_46_49333;
  wire seg_16_4_sp4_h_l_40_49460;
  wire seg_16_5_local_g1_2_64814;
  wire seg_16_5_local_g1_6_64818;
  wire seg_16_5_local_g2_0_64820;
  wire seg_16_5_local_g2_7_64827;
  wire seg_16_5_local_g3_1_64829;
  wire seg_16_5_local_g3_2_64830;
  wire seg_16_5_local_g3_3_64831;
  wire seg_16_5_local_g3_6_64834;
  wire seg_16_5_lutff_2_out_60934;
  wire seg_16_5_lutff_3_out_60935;
  wire seg_16_5_lutff_4_out_60936;
  wire seg_16_5_lutff_5_out_60937;
  wire seg_16_5_lutff_6_out_60938;
  wire seg_16_5_lutff_7_out_60939;
  wire seg_16_5_neigh_op_rgt_0_64763;
  wire seg_16_5_neigh_op_rgt_1_64764;
  wire seg_16_5_neigh_op_rgt_2_64765;
  wire seg_16_5_neigh_op_rgt_3_64766;
  wire seg_16_5_neigh_op_rgt_6_64769;
  wire seg_16_5_neigh_op_rgt_7_64770;
  wire seg_16_5_sp4_h_r_18_61076;
  wire seg_16_5_sp4_v_b_22_60843;
  wire seg_16_6_local_g2_0_64943;
  wire seg_16_6_lutff_0_out_61055;
  wire seg_16_6_neigh_op_rgt_0_64886;
  wire seg_16_6_sp4_h_l_36_49700;
  wire seg_16_6_sp4_h_l_41_49705;
  wire seg_16_6_sp4_h_l_42_49708;
  wire seg_16_6_sp4_h_r_6_65029;
  wire seg_16_6_sp4_v_b_6_60840;
  wire seg_16_7_sp4_v_b_8_60965;
  wire seg_16_8_sp4_v_b_5_61083;
  wire seg_16_9_glb_netwk_0_5;
  wire seg_16_9_local_g0_2_65298;
  wire seg_16_9_local_g0_6_65302;
  wire seg_16_9_local_g1_0_65304;
  wire seg_16_9_local_g1_3_65307;
  wire seg_16_9_local_g1_4_65308;
  wire seg_16_9_local_g2_3_65315;
  wire seg_16_9_local_g2_6_65318;
  wire seg_16_9_local_g3_1_65321;
  wire seg_16_9_lutff_2_out_61426;
  wire seg_16_9_lutff_3_out_61427;
  wire seg_16_9_lutff_4_out_61428;
  wire seg_16_9_lutff_5_out_61429;
  wire seg_16_9_lutff_6_out_61430;
  wire seg_16_9_sp12_v_b_14_64773;
  wire seg_16_9_sp4_r_v_b_14_65158;
  wire seg_16_9_sp4_r_v_b_17_65161;
  wire seg_16_9_sp4_v_b_0_61203;
  wire seg_16_9_sp4_v_b_19_61332;
  wire seg_16_9_sp4_v_b_36_61571;
  wire seg_16_9_sp4_v_b_44_61579;
  wire seg_16_9_sp4_v_b_4_61207;
  wire seg_17_0_glb_netwk_0_5;
  wire seg_17_0_local_g1_3_68056;
  wire seg_17_0_local_g1_5_68058;
  wire seg_17_0_span12_vert_16_68077;
  wire seg_17_0_span4_horz_r_0_68093;
  wire seg_17_0_span4_horz_r_11_60434;
  wire seg_17_0_span4_vert_16_64390;
  wire seg_17_0_span4_vert_18_64392;
  wire seg_17_0_span4_vert_21_64396;
  wire seg_17_10_sp4_h_l_36_54023;
  wire seg_17_10_sp4_h_l_37_54022;
  wire seg_17_10_sp4_h_r_10_69346;
  wire seg_17_10_sp4_h_r_11_69347;
  wire seg_17_11_sp4_v_b_10_65290;
  wire seg_17_12_glb_netwk_0_5;
  wire seg_17_12_local_g0_7_69503;
  wire seg_17_12_local_g3_5_69525;
  wire seg_17_12_sp4_h_l_37_54268;
  wire seg_17_12_sp4_h_r_18_65768;
  wire seg_17_12_sp4_h_r_3_69595;
  wire seg_17_12_sp4_v_b_15_65528;
  wire seg_17_12_sp4_v_b_29_65652;
  wire seg_17_12_sp4_v_b_3_65404;
  wire seg_17_12_sp4_v_t_39_65897;
  wire seg_17_13_glb_netwk_0_5;
  wire seg_17_13_glb_netwk_5_10;
  wire seg_17_13_glb_netwk_6_11;
  wire seg_17_13_local_g0_0_69619;
  wire seg_17_13_local_g0_4_69623;
  wire seg_17_13_local_g1_0_69627;
  wire seg_17_13_local_g1_2_69629;
  wire seg_17_13_local_g1_3_69630;
  wire seg_17_13_lutff_3_out_65750;
  wire seg_17_13_neigh_op_lft_0_61916;
  wire seg_17_13_neigh_op_lft_3_61919;
  wire seg_17_13_sp4_h_l_40_54398;
  wire seg_17_13_sp4_h_r_0_69713;
  wire seg_17_13_sp4_h_r_20_65893;
  wire seg_17_13_sp4_r_v_b_29_69606;
  wire seg_17_13_sp4_v_b_18_65654;
  wire seg_17_13_sp4_v_t_43_66024;
  wire seg_17_14_glb_netwk_0_5;
  wire seg_17_14_local_g0_0_69742;
  wire seg_17_14_local_g0_5_69747;
  wire seg_17_14_local_g0_7_69749;
  wire seg_17_14_local_g1_0_69750;
  wire seg_17_14_local_g1_3_69753;
  wire seg_17_14_local_g1_4_69754;
  wire seg_17_14_local_g1_6_69756;
  wire seg_17_14_local_g2_2_69760;
  wire seg_17_14_local_g2_5_69763;
  wire seg_17_14_lutff_0_out_65870;
  wire seg_17_14_lutff_2_out_65872;
  wire seg_17_14_lutff_3_out_65873;
  wire seg_17_14_lutff_4_out_65874;
  wire seg_17_14_lutff_5_out_65875;
  wire seg_17_14_lutff_7_out_65877;
  wire seg_17_14_neigh_op_top_0_65993;
  wire seg_17_14_sp4_h_l_37_54514;
  wire seg_17_14_sp4_h_l_38_54519;
  wire seg_17_14_sp4_h_l_44_54525;
  wire seg_17_14_sp4_h_r_0_69836;
  wire seg_17_14_sp4_h_r_13_66005;
  wire seg_17_14_sp4_h_r_20_66016;
  wire seg_17_14_sp4_h_r_26_62178;
  wire seg_17_14_sp4_h_r_3_69841;
  wire seg_17_14_sp4_h_r_6_69844;
  wire seg_17_14_sp4_h_r_7_69845;
  wire seg_17_14_sp4_r_v_b_27_69727;
  wire seg_17_14_sp4_v_b_0_65649;
  wire seg_17_14_sp4_v_b_10_65659;
  wire seg_17_14_sp4_v_b_11_65658;
  wire seg_17_14_sp4_v_b_23_65782;
  wire seg_17_14_sp4_v_b_5_65652;
  wire seg_17_15_glb_netwk_0_5;
  wire seg_17_15_glb_netwk_5_10;
  wire seg_17_15_glb_netwk_6_11;
  wire seg_17_15_local_g0_0_69865;
  wire seg_17_15_local_g0_2_69867;
  wire seg_17_15_local_g1_0_69873;
  wire seg_17_15_local_g1_2_69875;
  wire seg_17_15_local_g1_4_69877;
  wire seg_17_15_local_g1_5_69878;
  wire seg_17_15_local_g1_6_69879;
  wire seg_17_15_local_g1_7_69880;
  wire seg_17_15_lutff_0_out_65993;
  wire seg_17_15_lutff_4_out_65997;
  wire seg_17_15_neigh_op_bot_0_65870;
  wire seg_17_15_sp4_h_l_37_54637;
  wire seg_17_15_sp4_h_r_16_66135;
  wire seg_17_15_sp4_h_r_18_66137;
  wire seg_17_15_sp4_h_r_6_69967;
  wire seg_17_15_sp4_r_v_b_26_69851;
  wire seg_17_15_sp4_r_v_b_31_69854;
  wire seg_17_15_sp4_r_v_b_5_69606;
  wire seg_17_15_sp4_v_b_14_65896;
  wire seg_17_16_glb_netwk_0_5;
  wire seg_17_16_local_g1_7_70003;
  wire seg_17_16_local_g3_2_70014;
  wire seg_17_16_local_g3_5_70017;
  wire seg_17_16_lutff_1_out_66117;
  wire seg_17_16_sp4_h_r_14_66256;
  wire seg_17_16_sp4_h_r_23_66253;
  wire seg_17_16_sp4_h_r_30_62428;
  wire seg_17_16_sp4_r_v_b_18_69854;
  wire seg_17_16_sp4_v_b_29_66144;
  wire seg_17_16_sp4_v_b_6_65901;
  wire seg_17_16_sp4_v_b_8_65903;
  wire seg_17_17_glb_netwk_0_5;
  wire seg_17_17_glb_netwk_5_10;
  wire seg_17_17_glb_netwk_6_11;
  wire seg_17_17_local_g0_1_70112;
  wire seg_17_17_local_g0_2_70113;
  wire seg_17_17_local_g1_1_70120;
  wire seg_17_17_local_g1_2_70121;
  wire seg_17_17_local_g1_4_70123;
  wire seg_17_17_local_g1_5_70124;
  wire seg_17_17_local_g2_1_70128;
  wire seg_17_17_local_g3_1_70136;
  wire seg_17_17_local_g3_2_70137;
  wire seg_17_17_local_g3_3_70138;
  wire seg_17_17_local_g3_5_70140;
  wire seg_17_17_lutff_0_out_66239;
  wire seg_17_17_lutff_2_out_66241;
  wire seg_17_17_neigh_op_bnl_1_62286;
  wire seg_17_17_neigh_op_bot_1_66117;
  wire seg_17_17_neigh_op_lft_1_62409;
  wire seg_17_17_neigh_op_top_2_66364;
  wire seg_17_17_sp4_h_l_37_54883;
  wire seg_17_17_sp4_h_l_40_54890;
  wire seg_17_17_sp4_h_l_44_54894;
  wire seg_17_17_sp4_h_r_10_70207;
  wire seg_17_17_sp4_h_r_14_66379;
  wire seg_17_17_sp4_h_r_18_66383;
  wire seg_17_17_sp4_h_r_29_62550;
  wire seg_17_17_sp4_h_r_2_70209;
  wire seg_17_17_sp4_h_r_35_62546;
  wire seg_17_17_sp4_r_v_b_29_70098;
  wire seg_17_17_sp4_r_v_b_9_69856;
  wire seg_17_17_sp4_v_b_12_66140;
  wire seg_17_17_sp4_v_t_42_66515;
  wire seg_17_18_glb_netwk_0_5;
  wire seg_17_18_local_g0_2_70236;
  wire seg_17_18_local_g0_5_70239;
  wire seg_17_18_local_g1_1_70243;
  wire seg_17_18_local_g1_3_70245;
  wire seg_17_18_local_g1_5_70247;
  wire seg_17_18_local_g1_6_70248;
  wire seg_17_18_local_g2_4_70254;
  wire seg_17_18_lutff_0_out_66362;
  wire seg_17_18_lutff_1_out_66363;
  wire seg_17_18_lutff_2_out_66364;
  wire seg_17_18_lutff_4_out_66366;
  wire seg_17_18_neigh_op_lft_2_62533;
  wire seg_17_18_neigh_op_top_6_66491;
  wire seg_17_18_sp12_h_r_4_62662;
  wire seg_17_18_sp4_h_l_38_55011;
  wire seg_17_18_sp4_h_l_40_55013;
  wire seg_17_18_sp4_h_r_12_66498;
  wire seg_17_18_sp4_h_r_14_66502;
  wire seg_17_18_sp4_h_r_22_66500;
  wire seg_17_18_sp4_h_r_36_58837;
  wire seg_17_18_sp4_h_r_3_70333;
  wire seg_17_18_sp4_h_r_44_58847;
  wire seg_17_18_sp4_h_r_5_70335;
  wire seg_17_18_sp4_r_v_b_1_69971;
  wire seg_17_18_sp4_r_v_b_45_70349;
  wire seg_17_18_sp4_v_b_21_66272;
  wire seg_17_18_sp4_v_b_44_66517;
  wire seg_17_18_sp4_v_b_8_66149;
  wire seg_17_19_glb_netwk_0_5;
  wire seg_17_19_local_g0_1_70358;
  wire seg_17_19_local_g0_5_70362;
  wire seg_17_19_local_g0_6_70363;
  wire seg_17_19_local_g1_0_70365;
  wire seg_17_19_local_g1_6_70371;
  wire seg_17_19_local_g2_1_70374;
  wire seg_17_19_local_g2_2_70375;
  wire seg_17_19_local_g2_3_70376;
  wire seg_17_19_local_g2_6_70379;
  wire seg_17_19_local_g3_1_70382;
  wire seg_17_19_local_g3_4_70385;
  wire seg_17_19_local_g3_7_70388;
  wire seg_17_19_lutff_1_out_66486;
  wire seg_17_19_lutff_5_out_66490;
  wire seg_17_19_lutff_6_out_66491;
  wire seg_17_19_lutff_7_out_66492;
  wire seg_17_19_neigh_op_lft_1_62655;
  wire seg_17_19_neigh_op_lft_6_62660;
  wire seg_17_19_neigh_op_tnl_3_62780;
  wire seg_17_19_neigh_op_top_0_66608;
  wire seg_17_19_sp4_h_l_39_55133;
  wire seg_17_19_sp4_h_l_42_55138;
  wire seg_17_19_sp4_h_l_43_55137;
  wire seg_17_19_sp4_h_l_45_55139;
  wire seg_17_19_sp4_h_r_24_62789;
  wire seg_17_19_sp4_h_r_30_62797;
  wire seg_17_19_sp4_h_r_44_58970;
  wire seg_17_19_sp4_h_r_6_70459;
  wire seg_17_19_sp4_h_r_8_70461;
  wire seg_17_19_sp4_r_v_b_29_70344;
  wire seg_17_19_sp4_v_b_34_66520;
  wire seg_17_19_sp4_v_b_41_66637;
  wire seg_17_20_glb_netwk_0_5;
  wire seg_17_20_glb_netwk_3_8;
  wire seg_17_20_local_g1_1_70489;
  wire seg_17_20_local_g1_5_70493;
  wire seg_17_20_local_g1_6_70494;
  wire seg_17_20_local_g2_1_70497;
  wire seg_17_20_local_g2_5_70501;
  wire seg_17_20_local_g2_6_70502;
  wire seg_17_20_local_g2_7_70503;
  wire seg_17_20_local_g3_3_70507;
  wire seg_17_20_local_g3_4_70508;
  wire seg_17_20_lutff_0_out_66608;
  wire seg_17_20_lutff_1_out_66609;
  wire seg_17_20_lutff_2_out_66610;
  wire seg_17_20_lutff_5_out_66613;
  wire seg_17_20_lutff_6_out_66614;
  wire seg_17_20_neigh_op_lft_5_62782;
  wire seg_17_20_neigh_op_top_6_66737;
  wire seg_17_20_sp4_h_l_46_55255;
  wire seg_17_20_sp4_h_r_17_66749;
  wire seg_17_20_sp4_h_r_25_62913;
  wire seg_17_20_sp4_h_r_39_59086;
  wire seg_17_20_sp4_v_b_18_66515;
  wire seg_17_20_sp4_v_b_28_66637;
  wire seg_17_20_sp4_v_b_43_66762;
  wire seg_17_20_sp4_v_b_6_66393;
  wire seg_17_21_glb_netwk_0_5;
  wire seg_17_21_local_g0_2_70605;
  wire seg_17_21_local_g0_3_70606;
  wire seg_17_21_local_g2_1_70620;
  wire seg_17_21_lutff_6_out_66737;
  wire seg_17_21_sp4_h_l_41_55381;
  wire seg_17_21_sp4_r_v_b_11_70350;
  wire seg_17_21_sp4_r_v_b_27_70588;
  wire seg_17_21_sp4_v_b_10_66520;
  wire seg_17_21_sp4_v_b_41_66883;
  wire seg_17_21_sp4_v_b_9_66517;
  wire seg_17_24_sp4_v_b_6_66885;
  wire seg_17_25_sp4_v_b_9_67009;
  wire seg_17_28_sp4_v_b_9_67378;
  wire seg_17_29_local_g2_1_71604;
  wire seg_17_29_local_g2_5_71608;
  wire seg_17_29_local_g2_6_71609;
  wire seg_17_29_local_g3_3_71614;
  wire seg_17_29_neigh_op_bnl_1_63762;
  wire seg_17_29_neigh_op_bnl_3_63764;
  wire seg_17_29_neigh_op_bnl_5_63766;
  wire seg_17_29_neigh_op_bnl_6_63767;
  wire seg_17_29_sp4_r_v_b_29_71574;
  wire seg_17_2_sp4_h_l_39_53042;
  wire seg_17_2_sp4_v_b_5_64390;
  wire seg_17_2_sp4_v_b_7_64392;
  wire seg_17_31_glb_netwk_0_5;
  wire seg_17_31_local_g0_5_71851;
  wire seg_17_31_local_g1_5_71859;
  wire seg_17_31_span4_horz_r_5_68032;
  wire seg_17_31_span4_vert_13_67863;
  wire seg_17_31_span4_vert_8_67748;
  wire seg_17_3_sp4_h_l_43_53169;
  wire seg_17_4_sp4_h_l_37_53284;
  wire seg_17_5_glb_netwk_0_5;
  wire seg_17_5_local_g0_3_68638;
  wire seg_17_5_local_g1_2_68645;
  wire seg_17_5_local_g1_3_68646;
  wire seg_17_5_local_g1_4_68647;
  wire seg_17_5_local_g1_5_68648;
  wire seg_17_5_local_g1_6_68649;
  wire seg_17_5_local_g1_7_68650;
  wire seg_17_5_local_g2_0_68651;
  wire seg_17_5_local_g2_4_68655;
  wire seg_17_5_local_g3_0_68659;
  wire seg_17_5_local_g3_3_68662;
  wire seg_17_5_local_g3_7_68666;
  wire seg_17_5_lutff_0_out_64763;
  wire seg_17_5_lutff_1_out_64764;
  wire seg_17_5_lutff_2_out_64765;
  wire seg_17_5_lutff_3_out_64766;
  wire seg_17_5_lutff_5_out_64768;
  wire seg_17_5_lutff_6_out_64769;
  wire seg_17_5_lutff_7_out_64770;
  wire seg_17_5_neigh_op_lft_2_60934;
  wire seg_17_5_neigh_op_lft_3_60935;
  wire seg_17_5_neigh_op_lft_4_60936;
  wire seg_17_5_neigh_op_lft_5_60937;
  wire seg_17_5_neigh_op_lft_6_60938;
  wire seg_17_5_neigh_op_lft_7_60939;
  wire seg_17_5_neigh_op_tnr_0_68717;
  wire seg_17_5_sp4_h_r_3_68734;
  wire seg_17_5_sp4_r_v_b_12_68495;
  wire seg_17_6_glb_netwk_0_5;
  wire seg_17_6_local_g0_0_68758;
  wire seg_17_6_local_g0_1_68759;
  wire seg_17_6_local_g0_6_68764;
  wire seg_17_6_local_g1_0_68766;
  wire seg_17_6_local_g1_2_68768;
  wire seg_17_6_local_g1_3_68769;
  wire seg_17_6_local_g1_5_68771;
  wire seg_17_6_local_g1_7_68773;
  wire seg_17_6_local_g2_0_68774;
  wire seg_17_6_local_g2_7_68781;
  wire seg_17_6_local_g3_0_68782;
  wire seg_17_6_local_g3_5_68787;
  wire seg_17_6_lutff_0_out_64886;
  wire seg_17_6_lutff_4_out_64890;
  wire seg_17_6_lutff_5_out_64891;
  wire seg_17_6_lutff_7_out_64893;
  wire seg_17_6_neigh_op_bnr_5_68599;
  wire seg_17_6_neigh_op_bot_1_64764;
  wire seg_17_6_neigh_op_bot_2_64765;
  wire seg_17_6_neigh_op_bot_6_64769;
  wire seg_17_6_neigh_op_bot_7_64770;
  wire seg_17_6_neigh_op_lft_0_61055;
  wire seg_17_6_neigh_op_rgt_0_68717;
  wire seg_17_6_neigh_op_rgt_7_68724;
  wire seg_17_6_sp4_h_l_46_53533;
  wire seg_17_6_sp4_h_r_29_61197;
  wire seg_17_6_sp4_v_b_19_64794;
  wire seg_17_6_sp4_v_b_3_64666;
  wire seg_17_6_sp4_v_b_8_64673;
  wire seg_17_7_sp4_h_r_1_68976;
  wire seg_17_8_sp4_v_b_0_64911;
  wire seg_17_9_glb_netwk_0_5;
  wire seg_17_9_glb_netwk_3_8;
  wire seg_17_9_local_g3_0_69151;
  wire seg_17_9_lutff_1_out_65256;
  wire seg_17_9_sp12_v_b_0_68077;
  wire seg_17_9_sp4_v_b_34_65290;
  wire seg_18_0_glb_netwk_0_5;
  wire seg_18_0_local_g0_2_71878;
  wire seg_18_0_local_g1_1_71885;
  wire seg_18_0_span4_horz_r_4_68093;
  wire seg_18_0_span4_vert_17_68222;
  wire seg_18_0_span4_vert_42_68250;
  wire seg_18_10_local_g0_3_73084;
  wire seg_18_10_local_g0_4_73085;
  wire seg_18_10_local_g1_1_73090;
  wire seg_18_10_local_g3_0_73105;
  wire seg_18_10_sp4_h_l_40_57859;
  wire seg_18_10_sp4_h_l_44_57863;
  wire seg_18_10_sp4_h_l_45_57862;
  wire seg_18_10_sp4_h_r_17_69350;
  wire seg_18_10_sp4_h_r_19_69352;
  wire seg_18_10_sp4_h_r_22_69347;
  wire seg_18_10_sp4_h_r_38_61687;
  wire seg_18_10_sp4_h_r_4_73181;
  wire seg_18_10_sp4_h_r_6_73183;
  wire seg_18_10_sp4_v_b_22_69120;
  wire seg_18_10_sp4_v_b_32_69242;
  wire seg_18_11_sp4_h_l_41_57981;
  wire seg_18_12_glb_netwk_0_5;
  wire seg_18_12_local_g0_3_73330;
  wire seg_18_12_local_g3_3_73354;
  wire seg_18_12_local_g3_4_73355;
  wire seg_18_12_sp4_h_r_12_69591;
  wire seg_18_12_sp4_h_r_30_65767;
  wire seg_18_12_sp4_h_r_6_73429;
  wire seg_18_12_sp4_r_v_b_19_73194;
  wire seg_18_12_sp4_v_b_19_69363;
  wire seg_18_12_sp4_v_b_44_69610;
  wire seg_18_13_glb_netwk_0_5;
  wire seg_18_13_local_g0_2_73452;
  wire seg_18_13_local_g0_3_73453;
  wire seg_18_13_local_g0_4_73454;
  wire seg_18_13_local_g1_3_73461;
  wire seg_18_13_local_g1_4_73462;
  wire seg_18_13_local_g2_1_73467;
  wire seg_18_13_local_g2_7_73473;
  wire seg_18_13_local_g3_1_73475;
  wire seg_18_13_local_g3_4_73478;
  wire seg_18_13_local_g3_5_73479;
  wire seg_18_13_local_g3_7_73481;
  wire seg_18_13_lutff_1_out_69579;
  wire seg_18_13_neigh_op_lft_3_65750;
  wire seg_18_13_neigh_op_top_4_69705;
  wire seg_18_13_sp12_h_r_4_65878;
  wire seg_18_13_sp4_h_l_36_58222;
  wire seg_18_13_sp4_h_l_39_58225;
  wire seg_18_13_sp4_h_l_42_58230;
  wire seg_18_13_sp4_h_l_43_58229;
  wire seg_18_13_sp4_h_l_45_58231;
  wire seg_18_13_sp4_h_l_47_58223;
  wire seg_18_13_sp4_h_r_0_73544;
  wire seg_18_13_sp4_h_r_10_73546;
  wire seg_18_13_sp4_h_r_11_73547;
  wire seg_18_13_sp4_h_r_12_69714;
  wire seg_18_13_sp4_h_r_14_69718;
  wire seg_18_13_sp4_h_r_22_69716;
  wire seg_18_13_sp4_h_r_26_65886;
  wire seg_18_13_sp4_h_r_29_65889;
  wire seg_18_13_sp4_h_r_39_62055;
  wire seg_18_13_sp4_h_r_41_62057;
  wire seg_18_13_sp4_h_r_47_62053;
  wire seg_18_13_sp4_h_r_4_73550;
  wire seg_18_13_sp4_h_r_8_73554;
  wire seg_18_13_sp4_r_v_b_17_73315;
  wire seg_18_13_sp4_r_v_b_20_73318;
  wire seg_18_14_glb_netwk_0_5;
  wire seg_18_14_glb_netwk_5_10;
  wire seg_18_14_glb_netwk_6_11;
  wire seg_18_14_local_g0_1_73574;
  wire seg_18_14_local_g0_2_73575;
  wire seg_18_14_local_g0_3_73576;
  wire seg_18_14_local_g0_7_73580;
  wire seg_18_14_local_g1_1_73582;
  wire seg_18_14_local_g1_2_73583;
  wire seg_18_14_local_g1_4_73585;
  wire seg_18_14_local_g1_7_73588;
  wire seg_18_14_local_g2_0_73589;
  wire seg_18_14_local_g2_1_73590;
  wire seg_18_14_local_g2_2_73591;
  wire seg_18_14_local_g2_3_73592;
  wire seg_18_14_local_g2_6_73595;
  wire seg_18_14_local_g2_7_73596;
  wire seg_18_14_local_g3_2_73599;
  wire seg_18_14_local_g3_5_73602;
  wire seg_18_14_local_g3_7_73604;
  wire seg_18_14_lutff_1_out_69702;
  wire seg_18_14_lutff_4_out_69705;
  wire seg_18_14_lutff_7_out_69708;
  wire seg_18_14_neigh_op_bnr_1_73410;
  wire seg_18_14_neigh_op_bnr_7_73416;
  wire seg_18_14_neigh_op_bot_1_69579;
  wire seg_18_14_neigh_op_lft_2_65872;
  wire seg_18_14_neigh_op_lft_3_65873;
  wire seg_18_14_neigh_op_lft_4_65874;
  wire seg_18_14_neigh_op_lft_7_65877;
  wire seg_18_14_neigh_op_tnr_2_73657;
  wire seg_18_14_neigh_op_tnr_5_73660;
  wire seg_18_14_sp4_h_l_36_58345;
  wire seg_18_14_sp4_h_l_37_58344;
  wire seg_18_14_sp4_h_l_38_58349;
  wire seg_18_14_sp4_h_l_41_58350;
  wire seg_18_14_sp4_h_l_42_58353;
  wire seg_18_14_sp4_h_r_0_73667;
  wire seg_18_14_sp4_h_r_10_73669;
  wire seg_18_14_sp4_h_r_18_69845;
  wire seg_18_14_sp4_h_r_20_69847;
  wire seg_18_14_sp4_h_r_35_66008;
  wire seg_18_14_sp4_h_r_6_73675;
  wire seg_18_14_sp4_r_v_b_10_73321;
  wire seg_18_14_sp4_r_v_b_38_73681;
  wire seg_18_14_sp4_r_v_b_8_73319;
  wire seg_18_14_sp4_v_b_39_69851;
  wire seg_18_14_sp4_v_b_5_69483;
  wire seg_18_15_glb_netwk_0_5;
  wire seg_18_15_local_g0_5_73701;
  wire seg_18_15_local_g2_1_73713;
  wire seg_18_15_local_g2_5_73717;
  wire seg_18_15_local_g3_2_73722;
  wire seg_18_15_local_g3_3_73723;
  wire seg_18_15_local_g3_4_73724;
  wire seg_18_15_local_g3_5_73725;
  wire seg_18_15_sp4_h_l_38_58472;
  wire seg_18_15_sp4_h_l_44_58478;
  wire seg_18_15_sp4_h_r_0_73790;
  wire seg_18_15_sp4_h_r_13_69959;
  wire seg_18_15_sp4_h_r_14_69964;
  wire seg_18_15_sp4_h_r_20_69970;
  wire seg_18_15_sp4_h_r_27_66133;
  wire seg_18_15_sp4_h_r_28_66134;
  wire seg_18_15_sp4_h_r_34_66130;
  wire seg_18_15_sp4_h_r_40_62304;
  wire seg_18_15_sp4_h_r_41_62303;
  wire seg_18_15_sp4_h_r_44_62308;
  wire seg_18_15_sp4_h_r_45_62307;
  wire seg_18_15_sp4_r_v_b_11_73443;
  wire seg_18_15_sp4_r_v_b_7_73439;
  wire seg_18_15_sp4_v_b_37_69972;
  wire seg_18_16_glb_netwk_0_5;
  wire seg_18_16_local_g3_2_73845;
  wire seg_18_16_local_g3_6_73849;
  wire seg_18_16_lutff_2_out_69949;
  wire seg_18_16_sp4_h_r_20_70093;
  wire seg_18_16_sp4_h_r_4_73919;
  wire seg_18_16_sp4_r_v_b_22_73689;
  wire seg_18_16_sp4_r_v_b_37_73926;
  wire seg_18_16_sp4_r_v_b_5_73560;
  wire seg_18_16_sp4_v_b_3_69727;
  wire seg_18_17_glb_netwk_0_5;
  wire seg_18_17_local_g0_4_73946;
  wire seg_18_17_local_g0_6_73948;
  wire seg_18_17_local_g1_0_73950;
  wire seg_18_17_local_g1_3_73953;
  wire seg_18_17_local_g1_5_73955;
  wire seg_18_17_local_g1_6_73956;
  wire seg_18_17_local_g2_4_73962;
  wire seg_18_17_local_g2_7_73965;
  wire seg_18_17_local_g3_3_73969;
  wire seg_18_17_local_g3_4_73970;
  wire seg_18_17_local_g3_5_73971;
  wire seg_18_17_neigh_op_lft_0_66239;
  wire seg_18_17_neigh_op_top_4_70197;
  wire seg_18_17_sp4_h_l_36_58714;
  wire seg_18_17_sp4_h_r_0_74036;
  wire seg_18_17_sp4_h_r_10_74038;
  wire seg_18_17_sp4_h_r_11_74039;
  wire seg_18_17_sp4_h_r_12_70206;
  wire seg_18_17_sp4_h_r_14_70210;
  wire seg_18_17_sp4_h_r_22_70208;
  wire seg_18_17_sp4_h_r_28_66380;
  wire seg_18_17_sp4_h_r_2_74040;
  wire seg_18_17_sp4_h_r_30_66382;
  wire seg_18_17_sp4_h_r_38_62548;
  wire seg_18_17_sp4_h_r_4_74042;
  wire seg_18_17_sp4_h_r_8_74046;
  wire seg_18_17_sp4_h_r_9_74047;
  wire seg_18_17_sp4_r_v_b_19_73809;
  wire seg_18_17_sp4_r_v_b_20_73810;
  wire seg_18_17_sp4_r_v_b_21_73811;
  wire seg_18_17_sp4_v_b_21_69980;
  wire seg_18_17_sp4_v_b_47_70228;
  wire seg_18_17_sp4_v_t_40_70344;
  wire seg_18_17_sp4_v_t_46_70350;
  wire seg_18_18_glb_netwk_0_5;
  wire seg_18_18_glb_netwk_5_10;
  wire seg_18_18_glb_netwk_6_11;
  wire seg_18_18_local_g0_0_74065;
  wire seg_18_18_local_g0_3_74068;
  wire seg_18_18_local_g0_5_74070;
  wire seg_18_18_local_g0_7_74072;
  wire seg_18_18_local_g1_1_74074;
  wire seg_18_18_local_g1_3_74076;
  wire seg_18_18_local_g1_4_74077;
  wire seg_18_18_local_g1_7_74080;
  wire seg_18_18_local_g2_1_74082;
  wire seg_18_18_local_g2_2_74083;
  wire seg_18_18_local_g2_3_74084;
  wire seg_18_18_local_g2_5_74086;
  wire seg_18_18_local_g3_2_74091;
  wire seg_18_18_local_g3_3_74092;
  wire seg_18_18_lutff_3_out_70196;
  wire seg_18_18_lutff_4_out_70197;
  wire seg_18_18_lutff_5_out_70198;
  wire seg_18_18_neigh_op_bnr_7_73908;
  wire seg_18_18_neigh_op_lft_0_66362;
  wire seg_18_18_neigh_op_lft_1_66363;
  wire seg_18_18_neigh_op_lft_4_66366;
  wire seg_18_18_neigh_op_rgt_1_74025;
  wire seg_18_18_neigh_op_rgt_2_74026;
  wire seg_18_18_neigh_op_rgt_5_74029;
  wire seg_18_18_neigh_op_top_7_70323;
  wire seg_18_18_sp12_h_r_3_70324;
  wire seg_18_18_sp4_h_l_36_58837;
  wire seg_18_18_sp4_h_l_45_58846;
  wire seg_18_18_sp4_h_r_12_70329;
  wire seg_18_18_sp4_h_r_19_70336;
  wire seg_18_18_sp4_h_r_27_66502;
  wire seg_18_18_sp4_h_r_30_66505;
  wire seg_18_18_sp4_h_r_4_74165;
  wire seg_18_18_sp4_r_v_b_10_73813;
  wire seg_18_19_glb_netwk_0_5;
  wire seg_18_19_glb_netwk_5_10;
  wire seg_18_19_local_g0_7_74195;
  wire seg_18_19_lutff_7_out_70323;
  wire seg_18_19_sp4_h_l_46_58962;
  wire seg_18_19_sp4_h_r_23_70453;
  wire seg_18_20_glb_netwk_0_5;
  wire seg_18_20_local_g1_1_74320;
  wire seg_18_20_neigh_op_lft_1_66609;
  wire seg_18_20_sp4_h_l_47_59084;
  wire seg_18_20_sp4_r_v_b_31_74300;
  wire seg_18_21_sp4_v_b_8_70349;
  wire seg_18_22_sp4_v_t_41_70960;
  wire seg_18_23_sp4_v_t_42_71084;
  wire seg_18_23_sp4_v_t_43_71085;
  wire seg_18_25_sp4_h_r_10_75022;
  wire seg_18_25_sp4_v_b_4_70837;
  wire seg_18_26_sp4_v_t_36_71447;
  wire seg_18_27_sp4_v_t_41_71575;
  wire seg_18_27_sp4_v_t_43_71577;
  wire seg_18_29_sp4_v_b_10_71335;
  wire seg_18_2_sp4_h_l_47_56870;
  wire seg_18_30_sp4_v_t_36_75655;
  wire seg_18_31_glb_netwk_0_5;
  wire seg_18_31_local_g0_2_75679;
  wire seg_18_31_local_g0_5_75682;
  wire seg_18_31_span4_vert_34_71823;
  wire seg_18_31_span4_vert_36_75655;
  wire seg_18_31_span4_vert_4_71575;
  wire seg_18_31_span4_vert_5_71574;
  wire seg_18_31_span4_vert_6_71577;
  wire seg_18_4_sp4_h_l_36_57115;
  wire seg_18_5_glb_netwk_0_5;
  wire seg_18_5_local_g0_0_72466;
  wire seg_18_5_local_g1_5_72479;
  wire seg_18_5_local_g2_2_72484;
  wire seg_18_5_local_g2_3_72485;
  wire seg_18_5_local_g3_5_72495;
  wire seg_18_5_local_g3_7_72497;
  wire seg_18_5_lutff_5_out_68599;
  wire seg_18_5_lutff_7_out_68601;
  wire seg_18_5_neigh_op_top_0_68717;
  wire seg_18_5_sp4_h_r_26_64902;
  wire seg_18_5_sp4_h_r_42_61076;
  wire seg_18_5_sp4_v_b_13_68496;
  wire seg_18_5_sp4_v_b_43_68748;
  wire seg_18_6_glb_netwk_0_5;
  wire seg_18_6_local_g0_4_72593;
  wire seg_18_6_local_g0_5_72594;
  wire seg_18_6_local_g0_7_72596;
  wire seg_18_6_local_g1_0_72597;
  wire seg_18_6_local_g1_3_72600;
  wire seg_18_6_local_g1_4_72601;
  wire seg_18_6_local_g1_5_72602;
  wire seg_18_6_local_g1_7_72604;
  wire seg_18_6_local_g2_0_72605;
  wire seg_18_6_local_g2_2_72607;
  wire seg_18_6_local_g2_5_72610;
  wire seg_18_6_local_g2_7_72612;
  wire seg_18_6_local_g3_0_72613;
  wire seg_18_6_local_g3_5_72618;
  wire seg_18_6_lutff_0_out_68717;
  wire seg_18_6_lutff_2_out_68719;
  wire seg_18_6_lutff_5_out_68722;
  wire seg_18_6_lutff_7_out_68724;
  wire seg_18_6_neigh_op_bnl_5_64768;
  wire seg_18_6_neigh_op_bot_5_68599;
  wire seg_18_6_neigh_op_lft_4_64890;
  wire seg_18_6_neigh_op_lft_5_64891;
  wire seg_18_6_neigh_op_lft_7_64893;
  wire seg_18_6_sp4_h_l_42_57369;
  wire seg_18_6_sp4_h_r_10_72685;
  wire seg_18_6_sp4_h_r_24_65021;
  wire seg_18_6_sp4_h_r_2_72687;
  wire seg_18_6_sp4_h_r_30_65029;
  wire seg_18_6_sp4_h_r_44_61201;
  wire seg_18_6_sp4_h_r_4_72689;
  wire seg_18_6_sp4_h_r_7_72692;
  wire seg_18_6_sp4_r_v_b_16_72453;
  wire seg_18_6_sp4_r_v_b_3_72328;
  wire seg_18_7_sp4_v_t_46_69120;
  wire seg_18_8_sp4_h_l_45_57616;
  wire seg_19_10_sp4_h_l_42_61691;
  wire seg_19_10_sp4_h_r_0_76795;
  wire seg_19_10_sp4_h_r_10_76797;
  wire seg_19_10_sp4_h_r_3_76800;
  wire seg_19_12_sp4_h_l_36_61929;
  wire seg_19_12_sp4_v_b_11_73074;
  wire seg_19_12_sp4_v_b_6_73071;
  wire seg_19_12_sp4_v_t_43_73563;
  wire seg_19_13_glb_netwk_0_5;
  wire seg_19_13_local_g0_0_77027;
  wire seg_19_13_local_g0_3_77030;
  wire seg_19_13_local_g0_4_77031;
  wire seg_19_13_local_g0_6_77033;
  wire seg_19_13_local_g0_7_77034;
  wire seg_19_13_local_g1_0_77035;
  wire seg_19_13_local_g1_1_77036;
  wire seg_19_13_local_g1_3_77038;
  wire seg_19_13_local_g1_4_77039;
  wire seg_19_13_local_g1_5_77040;
  wire seg_19_13_local_g1_7_77042;
  wire seg_19_13_local_g2_1_77044;
  wire seg_19_13_local_g2_5_77048;
  wire seg_19_13_local_g2_6_77049;
  wire seg_19_13_local_g2_7_77050;
  wire seg_19_13_local_g3_3_77054;
  wire seg_19_13_local_g3_5_77056;
  wire seg_19_13_local_g3_6_77057;
  wire seg_19_13_ram_RDATA_10_73414;
  wire seg_19_13_ram_RDATA_12_73412;
  wire seg_19_13_ram_RDATA_13_73411;
  wire seg_19_13_ram_RDATA_14_73410;
  wire seg_19_13_ram_RDATA_8_73416;
  wire seg_19_13_sp4_h_l_37_62051;
  wire seg_19_13_sp4_h_l_41_62057;
  wire seg_19_13_sp4_h_l_46_62054;
  wire seg_19_13_sp4_h_l_47_62053;
  wire seg_19_13_sp4_h_r_0_77101;
  wire seg_19_13_sp4_h_r_11_77104;
  wire seg_19_13_sp4_h_r_14_73549;
  wire seg_19_13_sp4_h_r_15_73548;
  wire seg_19_13_sp4_h_r_16_73551;
  wire seg_19_13_sp4_h_r_19_73552;
  wire seg_19_13_sp4_h_r_20_73555;
  wire seg_19_13_sp4_h_r_24_69713;
  wire seg_19_13_sp4_h_r_30_69721;
  wire seg_19_13_sp4_h_r_38_65887;
  wire seg_19_13_sp4_h_r_41_65888;
  wire seg_19_13_sp4_h_r_44_65893;
  wire seg_19_13_sp4_h_r_47_65884;
  wire seg_19_13_sp4_h_r_4_77107;
  wire seg_19_13_sp4_h_r_5_77108;
  wire seg_19_13_sp4_h_r_8_77111;
  wire seg_19_13_sp4_h_r_9_77112;
  wire seg_19_13_sp4_r_v_b_19_76916;
  wire seg_19_13_sp4_r_v_b_21_76918;
  wire seg_19_13_sp4_v_b_37_73557;
  wire seg_19_13_sp4_v_b_7_73193;
  wire seg_19_13_sp4_v_t_41_73684;
  wire seg_19_14_glb_netwk_0_5;
  wire seg_19_14_local_g0_0_77129;
  wire seg_19_14_local_g0_1_77130;
  wire seg_19_14_local_g0_2_77131;
  wire seg_19_14_local_g0_3_77132;
  wire seg_19_14_local_g0_4_77133;
  wire seg_19_14_local_g0_5_77134;
  wire seg_19_14_local_g0_6_77135;
  wire seg_19_14_local_g1_0_77137;
  wire seg_19_14_local_g1_4_77141;
  wire seg_19_14_local_g1_5_77142;
  wire seg_19_14_local_g2_2_77147;
  wire seg_19_14_local_g2_5_77150;
  wire seg_19_14_local_g2_6_77151;
  wire seg_19_14_local_g2_7_77152;
  wire seg_19_14_local_g3_3_77156;
  wire seg_19_14_local_g3_4_77157;
  wire seg_19_14_local_g3_5_77158;
  wire seg_19_14_local_g3_7_77160;
  wire seg_19_14_ram_RDATA_1_73538;
  wire seg_19_14_ram_RDATA_2_73537;
  wire seg_19_14_ram_RDATA_5_73534;
  wire seg_19_14_sp4_h_l_36_62175;
  wire seg_19_14_sp4_h_l_37_62174;
  wire seg_19_14_sp4_h_l_44_62185;
  wire seg_19_14_sp4_h_l_45_62184;
  wire seg_19_14_sp4_h_r_16_73674;
  wire seg_19_14_sp4_h_r_17_73673;
  wire seg_19_14_sp4_h_r_20_73678;
  wire seg_19_14_sp4_h_r_29_69843;
  wire seg_19_14_sp4_h_r_39_66009;
  wire seg_19_14_sp4_h_r_3_77208;
  wire seg_19_14_sp4_h_r_4_77209;
  wire seg_19_14_sp4_h_r_5_77210;
  wire seg_19_14_sp4_h_r_8_77213;
  wire seg_19_14_sp4_r_v_b_0_76910;
  wire seg_19_14_sp4_r_v_b_26_77116;
  wire seg_19_14_sp4_r_v_b_30_77120;
  wire seg_19_14_sp4_r_v_b_32_77122;
  wire seg_19_14_sp4_r_v_b_34_77124;
  wire seg_19_14_sp4_r_v_b_38_77217;
  wire seg_19_14_sp4_r_v_b_3_76911;
  wire seg_19_14_sp4_r_v_b_41_77220;
  wire seg_19_14_sp4_r_v_b_44_77223;
  wire seg_19_14_sp4_r_v_b_47_77226;
  wire seg_19_14_sp4_r_v_b_5_76913;
  wire seg_19_14_sp4_r_v_b_7_76915;
  wire seg_19_14_sp4_v_b_10_73321;
  wire seg_19_14_sp4_v_b_29_73560;
  wire seg_19_14_sp4_v_b_35_73566;
  wire seg_19_14_sp4_v_b_47_73690;
  wire seg_19_14_sp4_v_b_6_73317;
  wire seg_19_15_glb_netwk_0_5;
  wire seg_19_15_local_g0_0_77231;
  wire seg_19_15_local_g0_1_77232;
  wire seg_19_15_local_g0_2_77233;
  wire seg_19_15_local_g0_3_77234;
  wire seg_19_15_local_g0_4_77235;
  wire seg_19_15_local_g0_5_77236;
  wire seg_19_15_local_g1_0_77239;
  wire seg_19_15_local_g1_1_77240;
  wire seg_19_15_local_g1_7_77246;
  wire seg_19_15_local_g2_0_77247;
  wire seg_19_15_local_g2_1_77248;
  wire seg_19_15_local_g2_4_77251;
  wire seg_19_15_local_g2_5_77252;
  wire seg_19_15_local_g2_7_77254;
  wire seg_19_15_local_g3_3_77258;
  wire seg_19_15_local_g3_5_77260;
  wire seg_19_15_local_g3_6_77261;
  wire seg_19_15_local_g3_7_77262;
  wire seg_19_15_ram_RDATA_10_73660;
  wire seg_19_15_ram_RDATA_12_73658;
  wire seg_19_15_ram_RDATA_13_73657;
  wire seg_19_15_ram_RDATA_14_73656;
  wire seg_19_15_ram_RDATA_15_73655;
  wire seg_19_15_sp4_h_l_36_62298;
  wire seg_19_15_sp4_h_l_40_62304;
  wire seg_19_15_sp4_h_l_41_62303;
  wire seg_19_15_sp4_h_l_44_62308;
  wire seg_19_15_sp4_h_l_45_62307;
  wire seg_19_15_sp4_h_r_0_77305;
  wire seg_19_15_sp4_h_r_14_73795;
  wire seg_19_15_sp4_h_r_16_73797;
  wire seg_19_15_sp4_h_r_17_73796;
  wire seg_19_15_sp4_h_r_19_73798;
  wire seg_19_15_sp4_h_r_23_73792;
  wire seg_19_15_sp4_h_r_38_66133;
  wire seg_19_15_sp4_h_r_39_66132;
  wire seg_19_15_sp4_h_r_40_66135;
  wire seg_19_15_sp4_h_r_43_66136;
  wire seg_19_15_sp4_h_r_45_66138;
  wire seg_19_15_sp4_h_r_9_77316;
  wire seg_19_15_sp4_r_v_b_13_77114;
  wire seg_19_15_sp4_v_b_11_73443;
  wire seg_19_15_sp4_v_b_13_73557;
  wire seg_19_15_sp4_v_b_18_73562;
  wire seg_19_15_sp4_v_b_20_73564;
  wire seg_19_15_sp4_v_b_25_73679;
  wire seg_19_15_sp4_v_b_28_73684;
  wire seg_19_15_sp4_v_b_29_73683;
  wire seg_19_15_sp4_v_b_31_73685;
  wire seg_19_15_sp4_v_b_32_73688;
  wire seg_19_15_sp4_v_b_7_73439;
  wire seg_19_16_glb_netwk_0_5;
  wire seg_19_16_local_g0_1_77334;
  wire seg_19_16_local_g0_6_77339;
  wire seg_19_16_local_g1_1_77342;
  wire seg_19_16_local_g1_2_77343;
  wire seg_19_16_local_g1_5_77346;
  wire seg_19_16_local_g2_0_77349;
  wire seg_19_16_local_g2_2_77351;
  wire seg_19_16_local_g2_4_77353;
  wire seg_19_16_local_g2_5_77354;
  wire seg_19_16_local_g2_7_77356;
  wire seg_19_16_local_g3_0_77357;
  wire seg_19_16_local_g3_1_77358;
  wire seg_19_16_local_g3_2_77359;
  wire seg_19_16_local_g3_3_77360;
  wire seg_19_16_local_g3_4_77361;
  wire seg_19_16_local_g3_5_77362;
  wire seg_19_16_local_g3_6_77363;
  wire seg_19_16_local_g3_7_77364;
  wire seg_19_16_neigh_op_lft_2_69949;
  wire seg_19_16_neigh_op_rgt_1_77264;
  wire seg_19_16_neigh_op_rgt_2_77265;
  wire seg_19_16_neigh_op_rgt_3_77266;
  wire seg_19_16_neigh_op_rgt_4_77267;
  wire seg_19_16_neigh_op_rgt_5_77268;
  wire seg_19_16_neigh_op_rgt_6_77269;
  wire seg_19_16_neigh_op_rgt_7_77270;
  wire seg_19_16_ram_RDATA_1_73784;
  wire seg_19_16_ram_RDATA_3_73782;
  wire seg_19_16_ram_RDATA_5_73780;
  wire seg_19_16_ram_RDATA_7_73778;
  wire seg_19_16_sp4_h_l_39_62424;
  wire seg_19_16_sp4_h_l_44_62431;
  wire seg_19_16_sp4_h_r_0_77407;
  wire seg_19_16_sp4_h_r_14_73918;
  wire seg_19_16_sp4_h_r_26_70086;
  wire seg_19_16_sp4_h_r_32_70092;
  wire seg_19_16_sp4_h_r_36_66252;
  wire seg_19_16_sp4_h_r_42_66260;
  wire seg_19_16_sp4_h_r_5_77414;
  wire seg_19_16_sp4_h_r_9_77418;
  wire seg_19_16_sp4_r_v_b_15_77218;
  wire seg_19_16_sp4_r_v_b_19_77222;
  wire seg_19_16_sp4_v_b_14_73681;
  wire seg_19_16_sp4_v_b_1_73556;
  wire seg_19_16_sp4_v_b_24_73803;
  wire seg_19_16_sp4_v_b_45_73934;
  wire seg_19_16_sp4_v_b_6_73563;
  wire seg_19_17_glb_netwk_0_5;
  wire seg_19_17_local_g0_0_77435;
  wire seg_19_17_local_g0_1_77436;
  wire seg_19_17_local_g0_2_77437;
  wire seg_19_17_local_g0_4_77439;
  wire seg_19_17_local_g0_5_77440;
  wire seg_19_17_local_g1_3_77446;
  wire seg_19_17_local_g1_4_77447;
  wire seg_19_17_local_g1_6_77449;
  wire seg_19_17_local_g1_7_77450;
  wire seg_19_17_local_g2_1_77452;
  wire seg_19_17_local_g2_2_77453;
  wire seg_19_17_local_g2_5_77456;
  wire seg_19_17_local_g2_6_77457;
  wire seg_19_17_local_g3_2_77461;
  wire seg_19_17_local_g3_3_77462;
  wire seg_19_17_local_g3_5_77464;
  wire seg_19_17_local_g3_7_77466;
  wire seg_19_17_ram_RDATA_10_73906;
  wire seg_19_17_ram_RDATA_11_73905;
  wire seg_19_17_ram_RDATA_12_73904;
  wire seg_19_17_ram_RDATA_8_73908;
  wire seg_19_17_sp4_h_l_38_62548;
  wire seg_19_17_sp4_h_l_41_62549;
  wire seg_19_17_sp4_h_r_0_77509;
  wire seg_19_17_sp4_h_r_11_77512;
  wire seg_19_17_sp4_h_r_12_74037;
  wire seg_19_17_sp4_h_r_16_74043;
  wire seg_19_17_sp4_h_r_18_74045;
  wire seg_19_17_sp4_h_r_1_77510;
  wire seg_19_17_sp4_h_r_26_70209;
  wire seg_19_17_sp4_h_r_28_70211;
  wire seg_19_17_sp4_h_r_2_77513;
  wire seg_19_17_sp4_h_r_30_70213;
  wire seg_19_17_sp4_h_r_31_70214;
  wire seg_19_17_sp4_h_r_33_70216;
  wire seg_19_17_sp4_h_r_34_70207;
  wire seg_19_17_sp4_h_r_3_77514;
  wire seg_19_17_sp4_h_r_4_77515;
  wire seg_19_17_sp4_h_r_5_77516;
  wire seg_19_17_sp4_h_r_7_77518;
  wire seg_19_17_sp4_r_v_b_19_77324;
  wire seg_19_17_sp4_r_v_b_21_77326;
  wire seg_19_17_sp4_r_v_b_5_77219;
  wire seg_19_17_sp4_v_b_14_73804;
  wire seg_19_17_sp4_v_b_37_74049;
  wire seg_19_17_sp4_v_t_40_74175;
  wire seg_19_18_glb_netwk_0_5;
  wire seg_19_18_local_g0_1_77538;
  wire seg_19_18_local_g0_2_77539;
  wire seg_19_18_local_g0_4_77541;
  wire seg_19_18_local_g0_5_77542;
  wire seg_19_18_local_g1_0_77545;
  wire seg_19_18_local_g1_3_77548;
  wire seg_19_18_local_g1_4_77549;
  wire seg_19_18_local_g1_5_77550;
  wire seg_19_18_local_g2_0_77553;
  wire seg_19_18_local_g2_2_77555;
  wire seg_19_18_local_g2_5_77558;
  wire seg_19_18_local_g2_6_77559;
  wire seg_19_18_local_g3_0_77561;
  wire seg_19_18_local_g3_1_77562;
  wire seg_19_18_local_g3_2_77563;
  wire seg_19_18_local_g3_3_77564;
  wire seg_19_18_local_g3_4_77565;
  wire seg_19_18_local_g3_7_77568;
  wire seg_19_18_ram_RDATA_0_74031;
  wire seg_19_18_ram_RDATA_1_74030;
  wire seg_19_18_ram_RDATA_2_74029;
  wire seg_19_18_ram_RDATA_4_74027;
  wire seg_19_18_ram_RDATA_5_74026;
  wire seg_19_18_ram_RDATA_6_74025;
  wire seg_19_18_ram_RDATA_7_74024;
  wire seg_19_18_sp4_h_l_37_62666;
  wire seg_19_18_sp4_h_l_38_62671;
  wire seg_19_18_sp4_h_l_45_62676;
  wire seg_19_18_sp4_h_r_0_77611;
  wire seg_19_18_sp4_h_r_12_74160;
  wire seg_19_18_sp4_h_r_27_70333;
  wire seg_19_18_sp4_h_r_31_70337;
  wire seg_19_18_sp4_h_r_32_70338;
  wire seg_19_18_sp4_h_r_41_66503;
  wire seg_19_18_sp4_h_r_45_66507;
  wire seg_19_18_sp4_r_v_b_10_77328;
  wire seg_19_18_sp4_r_v_b_14_77421;
  wire seg_19_18_sp4_r_v_b_16_77423;
  wire seg_19_18_sp4_r_v_b_18_77425;
  wire seg_19_18_sp4_r_v_b_20_77427;
  wire seg_19_18_sp4_r_v_b_26_77524;
  wire seg_19_18_sp4_r_v_b_29_77525;
  wire seg_19_18_sp4_r_v_b_34_77532;
  wire seg_19_18_sp4_r_v_b_4_77322;
  wire seg_19_18_sp4_v_b_13_73926;
  wire seg_19_18_sp4_v_b_19_73932;
  wire seg_19_18_sp4_v_b_40_74175;
  wire seg_19_18_sp4_v_t_42_74300;
  wire seg_19_19_sp4_h_l_37_62789;
  wire seg_19_25_sp12_h_r_22_36709;
  wire seg_19_4_sp4_h_l_47_60946;
  wire seg_19_6_sp4_h_l_44_61201;
  wire seg_19_6_sp4_h_r_2_76391;
  wire seg_19_7_sp4_h_r_5_76496;
  wire seg_19_8_sp4_v_b_3_72574;
  wire seg_20_10_glb_netwk_0_5;
  wire seg_20_10_local_g0_2_80114;
  wire seg_20_10_local_g0_5_80117;
  wire seg_20_10_local_g0_7_80119;
  wire seg_20_10_local_g1_1_80121;
  wire seg_20_10_local_g1_2_80122;
  wire seg_20_10_local_g1_3_80123;
  wire seg_20_10_local_g1_5_80125;
  wire seg_20_10_local_g2_1_80129;
  wire seg_20_10_local_g2_4_80132;
  wire seg_20_10_local_g3_0_80136;
  wire seg_20_10_local_g3_1_80137;
  wire seg_20_10_local_g3_3_80139;
  wire seg_20_10_local_g3_4_80140;
  wire seg_20_10_lutff_0_out_76651;
  wire seg_20_10_lutff_3_out_76654;
  wire seg_20_10_lutff_7_out_76658;
  wire seg_20_10_neigh_op_bot_1_76550;
  wire seg_20_10_neigh_op_bot_5_76554;
  wire seg_20_10_neigh_op_rgt_1_80072;
  wire seg_20_10_neigh_op_rgt_4_80075;
  wire seg_20_10_sp12_v_b_14_79589;
  wire seg_20_10_sp4_h_r_0_80206;
  wire seg_20_10_sp4_h_r_10_80208;
  wire seg_20_10_sp4_h_r_14_76800;
  wire seg_20_10_sp4_h_r_18_76804;
  wire seg_20_10_sp4_h_r_35_73178;
  wire seg_20_10_sp4_h_r_41_69350;
  wire seg_20_10_sp4_h_r_7_80215;
  wire seg_20_10_sp4_r_v_b_15_79975;
  wire seg_20_10_sp4_r_v_b_31_80101;
  wire seg_20_10_sp4_r_v_b_47_80229;
  wire seg_20_10_sp4_v_b_3_76503;
  wire seg_20_10_sp4_v_b_46_76817;
  wire seg_20_10_sp4_v_b_5_76505;
  wire seg_20_10_sp4_v_b_6_76508;
  wire seg_20_10_sp4_v_b_8_76510;
  wire seg_20_10_sp4_v_b_9_76509;
  wire seg_20_11_glb_netwk_0_5;
  wire seg_20_11_local_g0_7_80242;
  wire seg_20_11_lutff_5_out_76758;
  wire seg_20_11_sp4_v_b_15_76708;
  wire seg_20_12_glb_netwk_0_5;
  wire seg_20_12_glb_netwk_5_10;
  wire seg_20_12_glb_netwk_6_11;
  wire seg_20_12_local_g0_1_80359;
  wire seg_20_12_local_g0_2_80360;
  wire seg_20_12_local_g0_6_80364;
  wire seg_20_12_local_g1_2_80368;
  wire seg_20_12_local_g1_3_80369;
  wire seg_20_12_local_g1_5_80371;
  wire seg_20_12_local_g1_6_80372;
  wire seg_20_12_local_g1_7_80373;
  wire seg_20_12_local_g2_1_80375;
  wire seg_20_12_local_g2_2_80376;
  wire seg_20_12_local_g2_3_80377;
  wire seg_20_12_local_g2_4_80378;
  wire seg_20_12_local_g2_5_80379;
  wire seg_20_12_local_g2_6_80380;
  wire seg_20_12_local_g2_7_80381;
  wire seg_20_12_local_g3_3_80385;
  wire seg_20_12_local_g3_6_80388;
  wire seg_20_12_local_g3_7_80389;
  wire seg_20_12_lutff_0_out_76855;
  wire seg_20_12_lutff_1_out_76856;
  wire seg_20_12_lutff_2_out_76857;
  wire seg_20_12_lutff_3_out_76858;
  wire seg_20_12_lutff_4_out_76859;
  wire seg_20_12_lutff_5_out_76860;
  wire seg_20_12_lutff_6_out_76861;
  wire seg_20_12_lutff_7_out_76862;
  wire seg_20_12_neigh_op_bot_5_76758;
  wire seg_20_12_neigh_op_rgt_7_80324;
  wire seg_20_12_neigh_op_tnl_3_73412;
  wire seg_20_12_sp4_h_l_37_65759;
  wire seg_20_12_sp4_h_l_39_65763;
  wire seg_20_12_sp4_h_l_40_65766;
  wire seg_20_12_sp4_h_l_42_65768;
  wire seg_20_12_sp4_h_l_43_65767;
  wire seg_20_12_sp4_h_r_22_77002;
  wire seg_20_12_sp4_h_r_2_80456;
  wire seg_20_12_sp4_h_r_30_73429;
  wire seg_20_12_sp4_h_r_36_69591;
  wire seg_20_12_sp4_h_r_6_80460;
  wire seg_20_12_sp4_r_v_b_10_80106;
  wire seg_20_12_sp4_r_v_b_25_80341;
  wire seg_20_12_sp4_v_b_15_76810;
  wire seg_20_12_sp4_v_b_1_76705;
  wire seg_20_12_sp4_v_b_27_76911;
  wire seg_20_12_sp4_v_b_31_76915;
  wire seg_20_12_sp4_v_b_8_76714;
  wire seg_20_12_sp4_v_t_36_77113;
  wire seg_20_13_glb_netwk_0_5;
  wire seg_20_13_glb_netwk_5_10;
  wire seg_20_13_glb_netwk_6_11;
  wire seg_20_13_local_g0_0_80481;
  wire seg_20_13_local_g0_1_80482;
  wire seg_20_13_local_g0_2_80483;
  wire seg_20_13_local_g0_4_80485;
  wire seg_20_13_local_g0_5_80486;
  wire seg_20_13_local_g1_0_80489;
  wire seg_20_13_local_g1_2_80491;
  wire seg_20_13_local_g1_3_80492;
  wire seg_20_13_local_g1_4_80493;
  wire seg_20_13_local_g1_5_80494;
  wire seg_20_13_local_g1_6_80495;
  wire seg_20_13_local_g2_2_80499;
  wire seg_20_13_local_g2_4_80501;
  wire seg_20_13_local_g2_5_80502;
  wire seg_20_13_local_g2_6_80503;
  wire seg_20_13_local_g3_2_80507;
  wire seg_20_13_local_g3_4_80509;
  wire seg_20_13_local_g3_5_80510;
  wire seg_20_13_local_g3_6_80511;
  wire seg_20_13_lutff_0_out_76957;
  wire seg_20_13_lutff_4_out_76961;
  wire seg_20_13_lutff_7_out_76964;
  wire seg_20_13_neigh_op_bot_4_76859;
  wire seg_20_13_neigh_op_lft_2_73411;
  wire seg_20_13_neigh_op_lft_5_73414;
  wire seg_20_13_neigh_op_tnl_2_73534;
  wire seg_20_13_neigh_op_tnl_5_73537;
  wire seg_20_13_neigh_op_tnl_6_73538;
  wire seg_20_13_neigh_op_top_1_77060;
  wire seg_20_13_neigh_op_top_2_77061;
  wire seg_20_13_neigh_op_top_4_77063;
  wire seg_20_13_neigh_op_top_6_77065;
  wire seg_20_13_sp12_h_r_8_65878;
  wire seg_20_13_sp4_h_l_39_65886;
  wire seg_20_13_sp4_h_r_28_73550;
  wire seg_20_13_sp4_h_r_34_73546;
  wire seg_20_13_sp4_h_r_36_69714;
  wire seg_20_13_sp4_h_r_38_69718;
  wire seg_20_13_sp4_h_r_42_69722;
  wire seg_20_13_sp4_r_v_b_12_80341;
  wire seg_20_13_sp4_r_v_b_5_80222;
  wire seg_20_13_sp4_v_b_11_76817;
  wire seg_20_13_sp4_v_b_22_76919;
  wire seg_20_13_sp4_v_b_28_77016;
  wire seg_20_13_sp4_v_b_37_77114;
  wire seg_20_13_sp4_v_b_42_77119;
  wire seg_20_13_sp4_v_b_8_76816;
  wire seg_20_13_sp4_v_t_40_77219;
  wire seg_20_13_sp4_v_t_41_77220;
  wire seg_20_13_sp4_v_t_43_77222;
  wire seg_20_13_sp4_v_t_47_77226;
  wire seg_20_14_glb_netwk_0_5;
  wire seg_20_14_local_g0_0_80604;
  wire seg_20_14_local_g0_1_80605;
  wire seg_20_14_local_g0_5_80609;
  wire seg_20_14_local_g0_7_80611;
  wire seg_20_14_local_g1_0_80612;
  wire seg_20_14_local_g1_1_80613;
  wire seg_20_14_local_g1_6_80618;
  wire seg_20_14_local_g1_7_80619;
  wire seg_20_14_local_g2_0_80620;
  wire seg_20_14_local_g2_2_80622;
  wire seg_20_14_local_g2_3_80623;
  wire seg_20_14_local_g2_4_80624;
  wire seg_20_14_local_g2_6_80626;
  wire seg_20_14_local_g3_0_80628;
  wire seg_20_14_local_g3_3_80631;
  wire seg_20_14_local_g3_7_80635;
  wire seg_20_14_lutff_0_out_77059;
  wire seg_20_14_lutff_1_out_77060;
  wire seg_20_14_lutff_2_out_77061;
  wire seg_20_14_lutff_3_out_77062;
  wire seg_20_14_lutff_4_out_77063;
  wire seg_20_14_lutff_5_out_77064;
  wire seg_20_14_lutff_6_out_77065;
  wire seg_20_14_lutff_7_out_77066;
  wire seg_20_14_neigh_op_bnr_7_80447;
  wire seg_20_14_neigh_op_bot_7_76964;
  wire seg_20_14_neigh_op_top_1_77162;
  wire seg_20_14_sp4_h_l_43_66013;
  wire seg_20_14_sp4_h_r_24_73667;
  wire seg_20_14_sp4_h_r_27_73672;
  wire seg_20_14_sp4_h_r_30_73675;
  wire seg_20_14_sp4_h_r_31_73676;
  wire seg_20_14_sp4_h_r_34_73669;
  wire seg_20_14_sp4_h_r_44_69847;
  wire seg_20_14_sp4_h_r_6_80706;
  wire seg_20_14_sp4_r_v_b_16_80468;
  wire seg_20_14_sp4_r_v_b_24_80588;
  wire seg_20_14_sp4_v_b_11_76919;
  wire seg_20_14_sp4_v_b_1_76909;
  wire seg_20_14_sp4_v_b_27_77115;
  wire seg_20_14_sp4_v_b_6_76916;
  wire seg_20_14_sp4_v_b_8_76918;
  wire seg_20_14_sp4_v_t_41_77322;
  wire seg_20_15_glb_netwk_0_5;
  wire seg_20_15_glb_netwk_5_10;
  wire seg_20_15_glb_netwk_6_11;
  wire seg_20_15_local_g0_0_80727;
  wire seg_20_15_local_g0_2_80729;
  wire seg_20_15_local_g0_4_80731;
  wire seg_20_15_local_g1_0_80735;
  wire seg_20_15_local_g1_1_80736;
  wire seg_20_15_local_g1_3_80738;
  wire seg_20_15_local_g1_4_80739;
  wire seg_20_15_local_g1_5_80740;
  wire seg_20_15_local_g1_6_80741;
  wire seg_20_15_local_g2_0_80743;
  wire seg_20_15_local_g2_1_80744;
  wire seg_20_15_local_g2_2_80745;
  wire seg_20_15_local_g2_4_80747;
  wire seg_20_15_local_g2_6_80749;
  wire seg_20_15_local_g3_0_80751;
  wire seg_20_15_local_g3_1_80752;
  wire seg_20_15_local_g3_2_80753;
  wire seg_20_15_local_g3_4_80755;
  wire seg_20_15_local_g3_6_80757;
  wire seg_20_15_lutff_0_out_77161;
  wire seg_20_15_lutff_1_out_77162;
  wire seg_20_15_lutff_2_out_77163;
  wire seg_20_15_lutff_3_out_77164;
  wire seg_20_15_lutff_4_out_77165;
  wire seg_20_15_lutff_5_out_77166;
  wire seg_20_15_neigh_op_lft_0_73655;
  wire seg_20_15_neigh_op_lft_1_73656;
  wire seg_20_15_neigh_op_lft_3_73658;
  wire seg_20_15_neigh_op_tnl_0_73778;
  wire seg_20_15_neigh_op_tnl_2_73780;
  wire seg_20_15_neigh_op_tnl_4_73782;
  wire seg_20_15_neigh_op_tnl_6_73784;
  wire seg_20_15_sp4_h_r_16_77312;
  wire seg_20_15_sp4_h_r_18_77314;
  wire seg_20_15_sp4_h_r_21_77315;
  wire seg_20_15_sp4_h_r_22_77308;
  wire seg_20_15_sp4_h_r_24_73790;
  wire seg_20_15_sp4_h_r_38_69964;
  wire seg_20_15_sp4_h_r_44_69970;
  wire seg_20_15_sp4_r_v_b_10_80475;
  wire seg_20_15_sp4_v_b_12_77113;
  wire seg_20_15_sp4_v_b_14_77115;
  wire seg_20_15_sp4_v_b_25_77215;
  wire seg_20_15_sp4_v_b_4_77016;
  wire seg_20_16_glb_netwk_0_5;
  wire seg_20_16_local_g0_5_80855;
  wire seg_20_16_local_g1_1_80859;
  wire seg_20_16_local_g1_4_80862;
  wire seg_20_16_local_g1_6_80864;
  wire seg_20_16_local_g2_2_80868;
  wire seg_20_16_local_g2_4_80870;
  wire seg_20_16_local_g2_5_80871;
  wire seg_20_16_local_g3_3_80877;
  wire seg_20_16_local_g3_7_80881;
  wire seg_20_16_lutff_1_out_77264;
  wire seg_20_16_lutff_2_out_77265;
  wire seg_20_16_lutff_3_out_77266;
  wire seg_20_16_lutff_4_out_77267;
  wire seg_20_16_lutff_5_out_77268;
  wire seg_20_16_lutff_6_out_77269;
  wire seg_20_16_lutff_7_out_77270;
  wire seg_20_16_sp4_h_r_28_73919;
  wire seg_20_16_sp4_h_r_4_80950;
  wire seg_20_16_sp4_r_v_b_27_80835;
  wire seg_20_16_sp4_r_v_b_31_80839;
  wire seg_20_16_sp4_v_b_10_77124;
  wire seg_20_16_sp4_v_b_11_77123;
  wire seg_20_16_sp4_v_b_14_77217;
  wire seg_20_16_sp4_v_b_20_77223;
  wire seg_20_16_sp4_v_b_28_77322;
  wire seg_20_16_sp4_v_b_2_77116;
  wire seg_20_16_sp4_v_b_34_77328;
  wire seg_20_16_sp4_v_b_38_77421;
  wire seg_20_16_sp4_v_b_40_77423;
  wire seg_20_16_sp4_v_b_5_77117;
  wire seg_20_16_sp4_v_b_6_77120;
  wire seg_20_16_sp4_v_b_8_77122;
  wire seg_20_16_sp4_v_b_9_77121;
  wire seg_20_17_glb_netwk_0_5;
  wire seg_20_17_glb_netwk_5_10;
  wire seg_20_17_glb_netwk_6_11;
  wire seg_20_17_local_g0_2_80975;
  wire seg_20_17_local_g0_3_80976;
  wire seg_20_17_local_g0_4_80977;
  wire seg_20_17_local_g0_5_80978;
  wire seg_20_17_local_g0_6_80979;
  wire seg_20_17_local_g0_7_80980;
  wire seg_20_17_local_g1_3_80984;
  wire seg_20_17_local_g1_4_80985;
  wire seg_20_17_local_g1_5_80986;
  wire seg_20_17_local_g1_6_80987;
  wire seg_20_17_local_g2_0_80989;
  wire seg_20_17_local_g2_1_80990;
  wire seg_20_17_local_g2_2_80991;
  wire seg_20_17_local_g2_3_80992;
  wire seg_20_17_local_g2_4_80993;
  wire seg_20_17_local_g2_6_80995;
  wire seg_20_17_local_g2_7_80996;
  wire seg_20_17_local_g3_0_80997;
  wire seg_20_17_local_g3_1_80998;
  wire seg_20_17_local_g3_4_81001;
  wire seg_20_17_local_g3_5_81002;
  wire seg_20_17_local_g3_6_81003;
  wire seg_20_17_lutff_1_out_77366;
  wire seg_20_17_lutff_2_out_77367;
  wire seg_20_17_lutff_3_out_77368;
  wire seg_20_17_lutff_5_out_77370;
  wire seg_20_17_lutff_6_out_77371;
  wire seg_20_17_lutff_7_out_77372;
  wire seg_20_17_neigh_op_bot_4_77267;
  wire seg_20_17_neigh_op_bot_5_77268;
  wire seg_20_17_neigh_op_lft_4_73905;
  wire seg_20_17_neigh_op_rgt_4_80936;
  wire seg_20_17_neigh_op_rgt_6_80938;
  wire seg_20_17_neigh_op_tnl_0_74024;
  wire seg_20_17_neigh_op_tnl_6_74030;
  wire seg_20_17_sp12_v_b_1_79589;
  wire seg_20_17_sp4_h_l_38_66379;
  wire seg_20_17_sp4_h_l_39_66378;
  wire seg_20_17_sp4_h_l_43_66382;
  wire seg_20_17_sp4_h_r_19_77517;
  wire seg_20_17_sp4_h_r_1_81068;
  wire seg_20_17_sp4_h_r_26_74040;
  wire seg_20_17_sp4_h_r_2_81071;
  wire seg_20_17_sp4_h_r_32_74046;
  wire seg_20_17_sp4_h_r_36_70206;
  wire seg_20_17_sp4_h_r_3_81072;
  wire seg_20_17_sp4_h_r_41_70211;
  wire seg_20_17_sp4_r_v_b_15_80836;
  wire seg_20_17_sp4_r_v_b_1_80710;
  wire seg_20_17_sp4_r_v_b_30_80963;
  wire seg_20_17_sp4_r_v_b_5_80714;
  wire seg_20_17_sp4_r_v_b_9_80718;
  wire seg_20_17_sp4_v_b_11_77225;
  wire seg_20_18_glb_netwk_0_5;
  wire seg_20_18_glb_netwk_5_10;
  wire seg_20_18_glb_netwk_6_11;
  wire seg_20_18_local_g0_2_81098;
  wire seg_20_18_local_g0_3_81099;
  wire seg_20_18_local_g0_6_81102;
  wire seg_20_18_local_g0_7_81103;
  wire seg_20_18_local_g1_1_81105;
  wire seg_20_18_local_g1_3_81107;
  wire seg_20_18_local_g1_6_81110;
  wire seg_20_18_local_g1_7_81111;
  wire seg_20_18_local_g2_0_81112;
  wire seg_20_18_local_g2_3_81115;
  wire seg_20_18_local_g2_7_81119;
  wire seg_20_18_local_g3_0_81120;
  wire seg_20_18_local_g3_5_81125;
  wire seg_20_18_lutff_1_out_77468;
  wire seg_20_18_lutff_3_out_77470;
  wire seg_20_18_lutff_4_out_77471;
  wire seg_20_18_lutff_7_out_77474;
  wire seg_20_18_neigh_op_bnl_3_73904;
  wire seg_20_18_neigh_op_bnl_5_73906;
  wire seg_20_18_neigh_op_bnr_6_80938;
  wire seg_20_18_neigh_op_lft_3_74027;
  wire seg_20_18_neigh_op_lft_7_74031;
  wire seg_20_18_neigh_op_top_6_77575;
  wire seg_20_18_neigh_op_top_7_77576;
  wire seg_20_18_sp4_h_l_37_66497;
  wire seg_20_18_sp4_h_l_43_66505;
  wire seg_20_18_sp4_h_l_46_66500;
  wire seg_20_18_sp4_h_r_11_81193;
  wire seg_20_18_sp4_h_r_18_77620;
  wire seg_20_18_sp4_h_r_9_81201;
  wire seg_20_18_sp4_r_v_b_16_80960;
  wire seg_20_18_sp4_r_v_b_27_81081;
  wire seg_20_18_sp4_r_v_b_8_80842;
  wire seg_20_19_glb_netwk_0_5;
  wire seg_20_19_local_g2_1_81236;
  wire seg_20_19_local_g2_5_81240;
  wire seg_20_19_lutff_6_out_77575;
  wire seg_20_19_lutff_7_out_77576;
  wire seg_20_19_sp4_h_l_38_66625;
  wire seg_20_19_sp4_h_l_42_66629;
  wire seg_20_19_sp4_h_r_41_70457;
  wire seg_20_19_sp4_h_r_45_70461;
  wire seg_20_2_sp4_v_t_43_76100;
  wire seg_20_4_sp4_h_l_40_64782;
  wire seg_20_5_sp4_v_t_45_76408;
  wire seg_20_6_glb_netwk_0_5;
  wire seg_20_6_local_g0_2_79622;
  wire seg_20_6_local_g0_4_79624;
  wire seg_20_6_local_g1_0_79628;
  wire seg_20_6_local_g1_2_79630;
  wire seg_20_6_local_g1_7_79635;
  wire seg_20_6_local_g2_2_79638;
  wire seg_20_6_local_g2_5_79641;
  wire seg_20_6_local_g3_2_79646;
  wire seg_20_6_local_g3_5_79649;
  wire seg_20_6_lutff_2_out_76245;
  wire seg_20_6_lutff_5_out_76248;
  wire seg_20_6_lutff_7_out_76250;
  wire seg_20_6_neigh_op_rgt_5_79584;
  wire seg_20_6_neigh_op_top_0_76345;
  wire seg_20_6_sp4_h_l_38_65026;
  wire seg_20_6_sp4_h_l_41_65027;
  wire seg_20_6_sp4_h_r_20_76398;
  wire seg_20_6_sp4_h_r_26_72687;
  wire seg_20_6_sp4_h_r_34_72685;
  wire seg_20_6_sp4_h_r_4_79720;
  wire seg_20_6_sp4_r_v_b_33_79611;
  wire seg_20_6_sp4_v_t_43_76508;
  wire seg_20_7_local_g1_5_79756;
  wire seg_20_7_local_g2_2_79761;
  wire seg_20_7_lutff_0_out_76345;
  wire seg_20_7_neigh_op_bnr_5_79584;
  wire seg_20_7_sp4_h_r_16_76496;
  wire seg_20_7_sp4_r_v_b_1_79480;
  wire seg_20_7_sp4_r_v_b_33_79734;
  wire seg_20_7_sp4_v_b_26_76402;
  wire seg_20_7_sp4_v_b_32_76408;
  wire seg_20_8_sp4_v_b_5_76301;
  wire seg_20_9_glb_netwk_0_5;
  wire seg_20_9_local_g0_2_79991;
  wire seg_20_9_local_g1_0_79997;
  wire seg_20_9_local_g1_3_80000;
  wire seg_20_9_local_g1_7_80004;
  wire seg_20_9_local_g3_1_80014;
  wire seg_20_9_lutff_1_out_76550;
  wire seg_20_9_lutff_5_out_76554;
  wire seg_20_9_neigh_op_top_0_76651;
  wire seg_20_9_neigh_op_top_3_76654;
  wire seg_20_9_sp4_r_v_b_19_79856;
  wire seg_20_9_sp4_r_v_b_33_79980;
  wire seg_20_9_sp4_r_v_b_7_79732;
  wire seg_20_9_sp4_v_b_2_76402;
  wire seg_21_10_glb_netwk_0_5;
  wire seg_21_10_local_g0_0_83943;
  wire seg_21_10_local_g0_2_83945;
  wire seg_21_10_local_g0_3_83946;
  wire seg_21_10_local_g0_4_83947;
  wire seg_21_10_local_g1_5_83956;
  wire seg_21_10_local_g2_4_83963;
  wire seg_21_10_local_g2_5_83964;
  wire seg_21_10_local_g3_0_83967;
  wire seg_21_10_local_g3_5_83972;
  wire seg_21_10_lutff_0_out_80071;
  wire seg_21_10_lutff_1_out_80072;
  wire seg_21_10_lutff_4_out_80075;
  wire seg_21_10_neigh_op_bnl_5_76554;
  wire seg_21_10_neigh_op_lft_0_76651;
  wire seg_21_10_neigh_op_lft_3_76654;
  wire seg_21_10_sp12_v_b_18_83666;
  wire seg_21_10_sp4_h_r_10_84039;
  wire seg_21_10_sp4_h_r_13_80206;
  wire seg_21_10_sp4_h_r_18_80215;
  wire seg_21_10_sp4_h_r_20_80217;
  wire seg_21_10_sp4_h_r_24_76795;
  wire seg_21_10_sp4_h_r_2_84041;
  wire seg_21_10_sp4_h_r_34_76797;
  wire seg_21_10_sp4_h_r_37_73175;
  wire seg_21_10_sp4_h_r_8_84047;
  wire seg_21_10_sp4_r_v_b_25_83926;
  wire seg_21_10_sp4_v_b_18_79978;
  wire seg_21_10_sp4_v_b_1_79849;
  wire seg_21_10_sp4_v_b_24_80096;
  wire seg_21_10_sp4_v_b_34_80106;
  wire seg_21_10_sp4_v_b_40_80222;
  wire seg_21_10_sp4_v_b_4_79854;
  wire seg_21_10_sp4_v_b_6_79856;
  wire seg_21_11_sp4_v_b_2_79975;
  wire seg_21_11_sp4_v_b_7_79978;
  wire seg_21_11_sp4_v_t_36_80464;
  wire seg_21_12_glb_netwk_0_5;
  wire seg_21_12_local_g0_0_84189;
  wire seg_21_12_local_g0_7_84196;
  wire seg_21_12_local_g1_0_84197;
  wire seg_21_12_local_g1_5_84202;
  wire seg_21_12_local_g1_7_84204;
  wire seg_21_12_local_g3_4_84217;
  wire seg_21_12_lutff_2_out_80319;
  wire seg_21_12_lutff_7_out_80324;
  wire seg_21_12_neigh_op_lft_0_76855;
  wire seg_21_12_neigh_op_lft_7_76862;
  wire seg_21_12_sp4_h_r_13_80452;
  wire seg_21_12_sp4_h_r_28_77005;
  wire seg_21_12_sp4_h_r_7_84292;
  wire seg_21_12_sp4_v_b_0_80096;
  wire seg_21_12_sp4_v_b_10_80106;
  wire seg_21_12_sp4_v_b_16_80222;
  wire seg_21_12_sp4_v_b_1_80095;
  wire seg_21_12_sp4_v_b_23_80229;
  wire seg_21_12_sp4_v_b_42_80470;
  wire seg_21_12_sp4_v_b_7_80101;
  wire seg_21_13_glb_netwk_0_5;
  wire seg_21_13_glb_netwk_5_10;
  wire seg_21_13_glb_netwk_6_11;
  wire seg_21_13_local_g0_1_84313;
  wire seg_21_13_local_g0_2_84314;
  wire seg_21_13_local_g0_4_84316;
  wire seg_21_13_local_g0_7_84319;
  wire seg_21_13_local_g1_1_84321;
  wire seg_21_13_local_g1_2_84322;
  wire seg_21_13_local_g1_4_84324;
  wire seg_21_13_local_g1_5_84325;
  wire seg_21_13_local_g1_6_84326;
  wire seg_21_13_local_g1_7_84327;
  wire seg_21_13_local_g2_0_84328;
  wire seg_21_13_local_g2_5_84333;
  wire seg_21_13_local_g2_6_84334;
  wire seg_21_13_local_g2_7_84335;
  wire seg_21_13_local_g3_2_84338;
  wire seg_21_13_local_g3_5_84341;
  wire seg_21_13_local_g3_6_84342;
  wire seg_21_13_local_g3_7_84343;
  wire seg_21_13_lutff_1_out_80441;
  wire seg_21_13_lutff_2_out_80442;
  wire seg_21_13_lutff_6_out_80446;
  wire seg_21_13_lutff_7_out_80447;
  wire seg_21_13_neigh_op_bot_2_80319;
  wire seg_21_13_neigh_op_lft_4_76961;
  wire seg_21_13_neigh_op_rgt_2_84273;
  wire seg_21_13_sp4_h_l_42_69722;
  wire seg_21_13_sp4_h_l_46_69716;
  wire seg_21_13_sp4_h_r_14_80580;
  wire seg_21_13_sp4_h_r_17_80581;
  wire seg_21_13_sp4_h_r_23_80577;
  wire seg_21_13_sp4_h_r_24_77101;
  wire seg_21_13_sp4_h_r_31_77110;
  wire seg_21_13_sp4_h_r_37_73544;
  wire seg_21_13_sp4_h_r_45_73554;
  wire seg_21_13_sp4_r_v_b_22_84182;
  wire seg_21_13_sp4_r_v_b_41_84423;
  wire seg_21_13_sp4_v_b_10_80229;
  wire seg_21_13_sp4_v_b_12_80341;
  wire seg_21_13_sp4_v_b_15_80344;
  wire seg_21_13_sp4_v_b_32_80473;
  wire seg_21_13_sp4_v_b_38_80589;
  wire seg_21_13_sp4_v_b_39_80590;
  wire seg_21_13_sp4_v_b_5_80222;
  wire seg_21_13_sp4_v_t_43_80717;
  wire seg_21_14_glb_netwk_0_5;
  wire seg_21_14_local_g0_1_84436;
  wire seg_21_14_local_g0_2_84437;
  wire seg_21_14_local_g0_3_84438;
  wire seg_21_14_local_g0_4_84439;
  wire seg_21_14_local_g0_6_84441;
  wire seg_21_14_local_g0_7_84442;
  wire seg_21_14_local_g1_0_84443;
  wire seg_21_14_local_g1_1_84444;
  wire seg_21_14_local_g1_2_84445;
  wire seg_21_14_local_g1_3_84446;
  wire seg_21_14_local_g1_4_84447;
  wire seg_21_14_local_g1_5_84448;
  wire seg_21_14_local_g1_7_84450;
  wire seg_21_14_local_g2_1_84452;
  wire seg_21_14_local_g2_2_84453;
  wire seg_21_14_local_g2_3_84454;
  wire seg_21_14_local_g2_4_84455;
  wire seg_21_14_local_g2_5_84456;
  wire seg_21_14_local_g2_7_84458;
  wire seg_21_14_local_g3_0_84459;
  wire seg_21_14_local_g3_3_84462;
  wire seg_21_14_local_g3_4_84463;
  wire seg_21_14_local_g3_6_84465;
  wire seg_21_14_local_g3_7_84466;
  wire seg_21_14_lutff_1_out_80564;
  wire seg_21_14_lutff_2_out_80565;
  wire seg_21_14_lutff_3_out_80566;
  wire seg_21_14_lutff_4_out_80567;
  wire seg_21_14_lutff_5_out_80568;
  wire seg_21_14_lutff_7_out_80570;
  wire seg_21_14_neigh_op_bnl_0_76957;
  wire seg_21_14_neigh_op_bot_2_80442;
  wire seg_21_14_neigh_op_lft_3_77062;
  wire seg_21_14_neigh_op_lft_7_77066;
  wire seg_21_14_neigh_op_top_0_80686;
  wire seg_21_14_neigh_op_top_1_80687;
  wire seg_21_14_neigh_op_top_5_80691;
  wire seg_21_14_neigh_op_top_7_80693;
  wire seg_21_14_sp12_v_b_11_83667;
  wire seg_21_14_sp4_h_r_3_84534;
  wire seg_21_14_sp4_r_v_b_47_84552;
  wire seg_21_14_sp4_v_b_12_80464;
  wire seg_21_14_sp4_v_b_14_80466;
  wire seg_21_14_sp4_v_b_18_80470;
  wire seg_21_14_sp4_v_b_2_80344;
  wire seg_21_14_sp4_v_b_30_80594;
  wire seg_21_14_sp4_v_b_32_80596;
  wire seg_21_14_sp4_v_b_36_80710;
  wire seg_21_14_sp4_v_b_44_80718;
  wire seg_21_14_sp4_v_b_4_80346;
  wire seg_21_14_sp4_v_b_8_80350;
  wire seg_21_14_sp4_v_b_9_80349;
  wire seg_21_14_sp4_v_t_36_80833;
  wire seg_21_14_sp4_v_t_47_80844;
  wire seg_21_15_glb_netwk_0_5;
  wire seg_21_15_local_g0_0_84558;
  wire seg_21_15_local_g0_2_84560;
  wire seg_21_15_local_g0_3_84561;
  wire seg_21_15_local_g0_4_84562;
  wire seg_21_15_local_g0_5_84563;
  wire seg_21_15_local_g0_6_84564;
  wire seg_21_15_local_g1_0_84566;
  wire seg_21_15_local_g1_1_84567;
  wire seg_21_15_local_g1_2_84568;
  wire seg_21_15_local_g1_3_84569;
  wire seg_21_15_local_g1_4_84570;
  wire seg_21_15_local_g1_5_84571;
  wire seg_21_15_local_g1_6_84572;
  wire seg_21_15_local_g1_7_84573;
  wire seg_21_15_local_g2_1_84575;
  wire seg_21_15_local_g2_4_84578;
  wire seg_21_15_local_g2_7_84581;
  wire seg_21_15_local_g3_0_84582;
  wire seg_21_15_local_g3_1_84583;
  wire seg_21_15_local_g3_2_84584;
  wire seg_21_15_local_g3_3_84585;
  wire seg_21_15_local_g3_4_84586;
  wire seg_21_15_local_g3_7_84589;
  wire seg_21_15_lutff_0_out_80686;
  wire seg_21_15_lutff_1_out_80687;
  wire seg_21_15_lutff_2_out_80688;
  wire seg_21_15_lutff_3_out_80689;
  wire seg_21_15_lutff_4_out_80690;
  wire seg_21_15_lutff_5_out_80691;
  wire seg_21_15_lutff_6_out_80692;
  wire seg_21_15_lutff_7_out_80693;
  wire seg_21_15_neigh_op_lft_0_77161;
  wire seg_21_15_neigh_op_lft_2_77163;
  wire seg_21_15_neigh_op_lft_3_77164;
  wire seg_21_15_neigh_op_lft_5_77166;
  wire seg_21_15_neigh_op_tnr_7_84647;
  wire seg_21_15_neigh_op_top_3_80812;
  wire seg_21_15_sp4_h_l_43_69967;
  wire seg_21_15_sp4_h_r_9_84663;
  wire seg_21_15_sp4_r_v_b_12_84418;
  wire seg_21_15_sp4_r_v_b_17_84423;
  wire seg_21_15_sp4_v_b_12_80587;
  wire seg_21_15_sp4_v_b_14_80589;
  wire seg_21_15_sp4_v_b_18_80593;
  wire seg_21_15_sp4_v_b_21_80596;
  wire seg_21_15_sp4_v_b_23_80598;
  wire seg_21_15_sp4_v_b_28_80715;
  wire seg_21_15_sp4_v_b_31_80716;
  wire seg_21_15_sp4_v_b_32_80719;
  wire seg_21_15_sp4_v_b_41_80838;
  wire seg_21_15_sp4_v_b_5_80468;
  wire seg_21_15_sp4_v_b_8_80473;
  wire seg_21_15_sp4_v_t_38_80958;
  wire seg_21_16_glb_netwk_0_5;
  wire seg_21_16_glb_netwk_5_10;
  wire seg_21_16_local_g0_1_84682;
  wire seg_21_16_local_g0_5_84686;
  wire seg_21_16_local_g1_5_84694;
  wire seg_21_16_local_g1_7_84696;
  wire seg_21_16_local_g2_1_84698;
  wire seg_21_16_local_g3_1_84706;
  wire seg_21_16_local_g3_6_84711;
  wire seg_21_16_lutff_3_out_80812;
  wire seg_21_16_lutff_4_out_80813;
  wire seg_21_16_lutff_6_out_80815;
  wire seg_21_16_neigh_op_tnl_1_77366;
  wire seg_21_16_neigh_op_top_5_80937;
  wire seg_21_16_sp4_h_l_39_70086;
  wire seg_21_16_sp4_h_l_44_70093;
  wire seg_21_16_sp4_h_r_24_77407;
  wire seg_21_16_sp4_r_v_b_33_84672;
  wire seg_21_16_sp4_v_b_13_80711;
  wire seg_21_16_sp4_v_b_1_80587;
  wire seg_21_16_sp4_v_b_23_80721;
  wire seg_21_16_sp4_v_t_38_81081;
  wire seg_21_17_glb_netwk_0_5;
  wire seg_21_17_local_g0_2_84806;
  wire seg_21_17_local_g0_4_84808;
  wire seg_21_17_local_g1_0_84812;
  wire seg_21_17_local_g1_1_84813;
  wire seg_21_17_local_g1_2_84814;
  wire seg_21_17_local_g1_3_84815;
  wire seg_21_17_local_g1_5_84817;
  wire seg_21_17_local_g2_1_84821;
  wire seg_21_17_local_g2_2_84822;
  wire seg_21_17_local_g2_4_84824;
  wire seg_21_17_local_g2_5_84825;
  wire seg_21_17_local_g2_6_84826;
  wire seg_21_17_local_g2_7_84827;
  wire seg_21_17_local_g3_1_84829;
  wire seg_21_17_local_g3_2_84830;
  wire seg_21_17_local_g3_3_84831;
  wire seg_21_17_local_g3_4_84832;
  wire seg_21_17_local_g3_5_84833;
  wire seg_21_17_local_g3_6_84834;
  wire seg_21_17_local_g3_7_84835;
  wire seg_21_17_lutff_0_out_80932;
  wire seg_21_17_lutff_1_out_80933;
  wire seg_21_17_lutff_2_out_80934;
  wire seg_21_17_lutff_3_out_80935;
  wire seg_21_17_lutff_4_out_80936;
  wire seg_21_17_lutff_5_out_80937;
  wire seg_21_17_lutff_6_out_80938;
  wire seg_21_17_lutff_7_out_80939;
  wire seg_21_17_neigh_op_bnl_1_77264;
  wire seg_21_17_neigh_op_bnl_2_77265;
  wire seg_21_17_neigh_op_bnl_3_77266;
  wire seg_21_17_neigh_op_bnl_6_77269;
  wire seg_21_17_neigh_op_bnl_7_77270;
  wire seg_21_17_neigh_op_bot_4_80813;
  wire seg_21_17_neigh_op_lft_2_77367;
  wire seg_21_17_neigh_op_rgt_2_84765;
  wire seg_21_17_neigh_op_rgt_5_84768;
  wire seg_21_17_neigh_op_rgt_6_84769;
  wire seg_21_17_sp4_h_l_36_70206;
  wire seg_21_17_sp4_h_l_37_70205;
  wire seg_21_17_sp4_h_r_11_84901;
  wire seg_21_17_sp4_h_r_12_81068;
  wire seg_21_17_sp4_h_r_1_84899;
  wire seg_21_17_sp4_h_r_37_74036;
  wire seg_21_17_sp4_h_r_3_84903;
  wire seg_21_17_sp4_h_r_41_74042;
  wire seg_21_17_sp4_h_r_44_74047;
  wire seg_21_17_sp4_h_r_7_84907;
  wire seg_21_17_sp4_r_v_b_12_84664;
  wire seg_21_17_sp4_r_v_b_13_84665;
  wire seg_21_17_sp4_v_b_12_80833;
  wire seg_21_17_sp4_v_b_44_81087;
  wire seg_21_18_glb_netwk_0_5;
  wire seg_21_18_glb_netwk_5_10;
  wire seg_21_18_local_g0_1_84928;
  wire seg_21_18_local_g0_2_84929;
  wire seg_21_18_local_g0_3_84930;
  wire seg_21_18_local_g0_4_84931;
  wire seg_21_18_local_g1_0_84935;
  wire seg_21_18_local_g1_1_84936;
  wire seg_21_18_local_g1_3_84938;
  wire seg_21_18_local_g1_4_84939;
  wire seg_21_18_local_g1_5_84940;
  wire seg_21_18_local_g1_6_84941;
  wire seg_21_18_local_g3_1_84952;
  wire seg_21_18_local_g3_2_84953;
  wire seg_21_18_local_g3_4_84955;
  wire seg_21_18_local_g3_6_84957;
  wire seg_21_18_lutff_1_out_81056;
  wire seg_21_18_lutff_3_out_81058;
  wire seg_21_18_lutff_4_out_81059;
  wire seg_21_18_lutff_6_out_81061;
  wire seg_21_18_neigh_op_lft_1_77468;
  wire seg_21_18_neigh_op_lft_3_77470;
  wire seg_21_18_neigh_op_lft_4_77471;
  wire seg_21_18_neigh_op_top_2_81180;
  wire seg_21_18_sp12_h_r_8_70324;
  wire seg_21_18_sp12_v_b_2_83666;
  wire seg_21_18_sp4_h_l_36_70329;
  wire seg_21_18_sp4_h_r_14_81195;
  wire seg_21_18_sp4_h_r_41_74165;
  wire seg_21_18_sp4_h_r_4_85027;
  wire seg_21_18_sp4_v_b_10_80844;
  wire seg_21_18_sp4_v_b_14_80958;
  wire seg_21_18_sp4_v_b_1_80833;
  wire seg_21_18_sp4_v_b_21_80965;
  wire seg_21_18_sp4_v_b_3_80835;
  wire seg_21_18_sp4_v_b_4_80838;
  wire seg_21_18_sp4_v_b_7_80839;
  wire seg_21_18_sp4_v_b_8_80842;
  wire seg_21_19_glb_netwk_0_5;
  wire seg_21_19_glb_netwk_5_10;
  wire seg_21_19_local_g1_6_85064;
  wire seg_21_19_lutff_2_out_81180;
  wire seg_21_19_sp4_h_l_47_70453;
  wire seg_21_19_sp4_h_r_6_85152;
  wire seg_21_19_sp4_v_b_6_80963;
  wire seg_21_5_sp4_v_t_44_79734;
  wire seg_21_6_local_g0_5_83456;
  wire seg_21_6_local_g1_1_83460;
  wire seg_21_6_local_g1_7_83466;
  wire seg_21_6_lutff_5_out_79584;
  wire seg_21_6_neigh_op_lft_5_76248;
  wire seg_21_6_neigh_op_lft_7_76250;
  wire seg_21_6_sp12_v_b_10_82776;
  wire seg_21_6_sp4_h_l_39_68856;
  wire seg_21_6_sp4_h_r_10_83547;
  wire seg_21_6_sp4_h_r_26_76391;
  wire seg_21_6_sp4_h_r_42_72692;
  wire seg_21_6_sp4_r_v_b_11_83198;
  wire seg_21_6_sp4_r_v_b_43_83564;
  wire seg_21_6_sp4_r_v_b_7_83194;
  wire seg_21_6_sp4_v_b_10_79368;
  wire seg_21_6_sp4_v_b_17_79485;
  wire seg_21_6_sp4_v_b_42_79732;
  wire seg_21_7_sp4_v_b_1_79480;
  wire seg_21_7_sp4_v_t_41_79977;
  wire seg_21_9_glb_netwk_0_5;
  wire seg_21_9_local_g0_2_83822;
  wire seg_21_9_local_g1_0_83828;
  wire seg_21_9_local_g1_5_83833;
  wire seg_21_9_local_g1_7_83835;
  wire seg_21_9_local_g2_7_83843;
  wire seg_21_9_local_g3_5_83849;
  wire seg_21_9_lutff_0_out_79948;
  wire seg_21_9_lutff_2_out_79950;
  wire seg_21_9_neigh_op_lft_5_76554;
  wire seg_21_9_sp12_v_b_20_83667;
  wire seg_21_9_sp12_v_b_5_82776;
  wire seg_21_9_sp4_h_r_0_83914;
  wire seg_21_9_sp4_h_r_20_80094;
  wire seg_21_9_sp4_h_r_28_76699;
  wire seg_21_9_sp4_r_v_b_15_83683;
  wire seg_21_9_sp4_v_b_15_79852;
  wire seg_21_9_sp4_v_b_36_80095;
  wire seg_21_9_sp4_v_b_7_79732;
  wire seg_22_0_local_g1_2_86579;
  wire seg_22_0_span4_vert_18_82916;
  wire seg_22_10_sp4_h_l_43_73183;
  wire seg_22_12_sp4_v_b_1_83926;
  wire seg_22_13_glb_netwk_0_5;
  wire seg_22_13_local_g1_1_88152;
  wire seg_22_13_local_g2_7_88166;
  wire seg_22_13_lutff_2_out_84273;
  wire seg_22_13_sp4_h_l_36_73545;
  wire seg_22_13_sp4_h_r_42_77110;
  wire seg_22_13_sp4_h_r_9_88248;
  wire seg_22_13_sp4_r_v_b_15_88006;
  wire seg_22_13_sp4_v_t_43_84548;
  wire seg_22_13_sp4_v_t_45_84550;
  wire seg_22_14_glb_netwk_0_5;
  wire seg_22_14_glb_netwk_5_10;
  wire seg_22_14_glb_netwk_6_11;
  wire seg_22_14_local_g0_4_88270;
  wire seg_22_14_local_g1_4_88278;
  wire seg_22_14_local_g1_5_88279;
  wire seg_22_14_neigh_op_top_4_84521;
  wire seg_22_14_sp4_h_l_40_73674;
  wire seg_22_14_sp4_h_r_38_77208;
  wire seg_22_14_sp4_h_r_5_88367;
  wire seg_22_14_sp4_v_b_20_84303;
  wire seg_22_14_sp4_v_b_6_84179;
  wire seg_22_14_sp4_v_t_37_84665;
  wire seg_22_15_glb_netwk_0_5;
  wire seg_22_15_local_g3_4_88417;
  wire seg_22_15_local_g3_6_88419;
  wire seg_22_15_lutff_4_out_84521;
  wire seg_22_15_sp4_h_l_38_73795;
  wire seg_22_15_sp4_h_r_44_77316;
  wire seg_22_15_sp4_r_v_b_37_88496;
  wire seg_22_15_sp4_v_b_36_84664;
  wire seg_22_15_sp4_v_b_38_84666;
  wire seg_22_15_sp4_v_t_41_84792;
  wire seg_22_15_sp4_v_t_47_84798;
  wire seg_22_16_glb_netwk_0_5;
  wire seg_22_16_glb_netwk_5_10;
  wire seg_22_16_glb_netwk_6_11;
  wire seg_22_16_local_g2_6_88534;
  wire seg_22_16_local_g3_3_88539;
  wire seg_22_16_lutff_7_out_84647;
  wire seg_22_16_neigh_op_tnl_6_80938;
  wire seg_22_16_sp4_r_v_b_19_88379;
  wire seg_22_17_local_g0_1_88636;
  wire seg_22_17_local_g0_3_88638;
  wire seg_22_17_local_g0_4_88639;
  wire seg_22_17_local_g0_5_88640;
  wire seg_22_17_local_g0_7_88642;
  wire seg_22_17_local_g1_3_88646;
  wire seg_22_17_local_g1_4_88647;
  wire seg_22_17_local_g1_7_88650;
  wire seg_22_17_local_g2_5_88656;
  wire seg_22_17_lutff_2_out_84765;
  wire seg_22_17_lutff_5_out_84768;
  wire seg_22_17_lutff_6_out_84769;
  wire seg_22_17_neigh_op_lft_3_80935;
  wire seg_22_17_neigh_op_lft_4_80936;
  wire seg_22_17_neigh_op_lft_5_80937;
  wire seg_22_17_neigh_op_lft_7_80939;
  wire seg_22_17_sp4_h_l_37_74036;
  wire seg_22_17_sp4_h_l_41_74042;
  wire seg_22_17_sp4_h_l_47_74038;
  wire seg_22_17_sp4_h_r_12_84899;
  wire seg_22_17_sp4_h_r_14_84903;
  wire seg_22_17_sp4_h_r_17_84904;
  wire seg_22_17_sp4_h_r_18_84907;
  wire seg_22_17_sp4_h_r_22_84901;
  wire seg_22_17_sp4_h_r_36_77510;
  wire seg_22_17_sp4_h_r_38_77514;
  wire seg_22_17_sp4_h_r_3_88734;
  wire seg_22_17_sp4_h_r_40_77516;
  wire seg_22_17_sp4_h_r_42_77518;
  wire seg_22_17_sp4_h_r_46_77512;
  wire seg_22_17_sp4_h_r_4_88735;
  wire seg_22_17_sp4_h_r_8_88739;
  wire seg_22_17_sp4_r_v_b_11_88382;
  wire seg_22_17_sp4_r_v_b_13_88496;
  wire seg_22_17_sp4_r_v_b_3_88374;
  wire seg_22_17_sp4_r_v_b_5_88376;
  wire seg_22_17_sp4_v_b_14_84666;
  wire seg_22_17_sp4_v_b_15_84667;
  wire seg_22_17_sp4_v_b_28_84792;
  wire seg_22_17_sp4_v_b_2_84544;
  wire seg_22_17_sp4_v_b_34_84798;
  wire seg_22_17_sp4_v_b_6_84548;
  wire seg_22_17_sp4_v_b_8_84550;
  wire seg_22_2_sp4_v_t_42_83194;
  wire seg_22_6_sp4_h_l_39_72687;
  wire seg_22_6_sp4_v_b_11_83198;
  wire seg_22_9_glb_netwk_0_5;
  wire seg_22_9_local_g0_1_87652;
  wire seg_22_9_local_g0_4_87655;
  wire seg_22_9_local_g2_2_87669;
  wire seg_22_9_lutff_1_out_83780;
  wire seg_22_9_sp4_h_r_12_83915;
  wire seg_22_9_sp4_r_v_b_10_87399;
  wire seg_22_9_sp4_v_b_6_83564;
  wire seg_23_13_sp4_v_t_38_88374;
  wire seg_23_13_sp4_v_t_40_88376;
  wire seg_23_13_sp4_v_t_46_88382;
  wire seg_23_14_sp4_h_l_45_77213;
  wire seg_23_17_sp4_h_l_37_77509;
  wire seg_23_6_sp4_v_t_38_87513;
  wire seg_23_9_glb_netwk_0_5;
  wire seg_23_9_local_g0_2_91484;
  wire seg_23_9_local_g1_1_91491;
  wire seg_23_9_local_g1_3_91493;
  wire seg_23_9_local_g1_5_91495;
  wire seg_23_9_local_g3_0_91506;
  wire seg_23_9_lutff_2_out_87612;
  wire seg_23_9_neigh_op_lft_1_83780;
  wire seg_23_9_sp4_h_l_41_76699;
  wire seg_23_9_sp4_h_r_13_87745;
  wire seg_23_9_sp4_h_r_24_83914;
  wire seg_23_9_sp4_r_v_b_3_91221;
  wire seg_23_9_sp4_v_b_14_87513;
  wire seg_24_9_sp4_h_l_44_80094;
  wire seg_2_19_local_g2_4_13545;
  wire seg_2_19_local_g3_2_13551;
  wire seg_2_19_local_g3_5_13554;
  wire seg_2_19_local_g3_6_13555;
  wire seg_2_19_neigh_op_rgt_4_13488;
  wire seg_2_19_neigh_op_rgt_5_13489;
  wire seg_2_19_neigh_op_rgt_6_13490;
  wire seg_2_19_neigh_op_tnr_2_13609;
  wire seg_2_19_sp4_h_r_0_13619;
  wire seg_2_8_glb_netwk_0_5;
  wire seg_2_8_local_g0_6_12178;
  wire seg_2_8_local_g0_7_12179;
  wire seg_2_8_local_g1_5_12185;
  wire seg_2_8_local_g2_3_12191;
  wire seg_2_8_local_g2_4_12192;
  wire seg_2_8_local_g3_2_12198;
  wire seg_2_8_local_g3_4_12200;
  wire seg_2_8_local_g3_5_12201;
  wire seg_2_8_lutff_2_out_7745;
  wire seg_2_8_lutff_3_out_7746;
  wire seg_2_8_lutff_4_out_7747;
  wire seg_2_8_lutff_5_out_7748;
  wire seg_2_8_lutff_6_out_7749;
  wire seg_2_8_neigh_op_bnr_7_12015;
  wire seg_2_8_neigh_op_rgt_4_12135;
  wire seg_2_8_sp4_h_r_46_1816;
  wire seg_2_8_sp4_r_v_b_15_12035;
  wire seg_2_8_sp4_r_v_b_5_11913;
  wire seg_3_13_glb_netwk_0_5;
  wire seg_3_13_local_g0_2_16620;
  wire seg_3_13_local_g1_2_16628;
  wire seg_3_13_local_g1_5_16631;
  wire seg_3_13_local_g1_6_16632;
  wire seg_3_13_local_g2_5_16639;
  wire seg_3_13_local_g3_3_16645;
  wire seg_3_13_local_g3_4_16646;
  wire seg_3_13_local_g3_5_16647;
  wire seg_3_13_lutff_2_out_12748;
  wire seg_3_13_lutff_3_out_12749;
  wire seg_3_13_lutff_4_out_12750;
  wire seg_3_13_lutff_5_out_12751;
  wire seg_3_13_lutff_6_out_12752;
  wire seg_3_13_neigh_op_rgt_5_16582;
  wire seg_3_13_neigh_op_top_2_12871;
  wire seg_3_13_sp12_v_b_14_16095;
  wire seg_3_13_sp4_h_r_14_12886;
  wire seg_3_13_sp4_h_r_46_2864;
  wire seg_3_13_sp4_r_v_b_5_16359;
  wire seg_3_14_glb_netwk_0_5;
  wire seg_3_14_local_g2_2_16759;
  wire seg_3_14_local_g3_3_16768;
  wire seg_3_14_local_g3_5_16770;
  wire seg_3_14_lutff_2_out_12871;
  wire seg_3_14_sp12_v_b_13_16095;
  wire seg_3_14_sp4_r_v_b_43_16854;
  wire seg_3_18_glb_netwk_0_5;
  wire seg_3_18_local_g0_4_17237;
  wire seg_3_18_local_g0_5_17238;
  wire seg_3_18_local_g0_6_17239;
  wire seg_3_18_local_g1_1_17242;
  wire seg_3_18_local_g2_2_17251;
  wire seg_3_18_local_g2_3_17252;
  wire seg_3_18_local_g2_7_17256;
  wire seg_3_18_local_g3_7_17264;
  wire seg_3_18_lutff_2_out_13363;
  wire seg_3_18_lutff_3_out_13364;
  wire seg_3_18_lutff_4_out_13365;
  wire seg_3_18_lutff_5_out_13366;
  wire seg_3_18_lutff_6_out_13367;
  wire seg_3_18_lutff_7_out_13368;
  wire seg_3_18_neigh_op_bnr_1_17070;
  wire seg_3_18_neigh_op_rgt_7_17199;
  wire seg_3_19_glb_netwk_0_5;
  wire seg_3_19_local_g0_1_17357;
  wire seg_3_19_local_g0_6_17362;
  wire seg_3_19_local_g1_0_17364;
  wire seg_3_19_local_g1_3_17367;
  wire seg_3_19_local_g2_4_17376;
  wire seg_3_19_local_g2_5_17377;
  wire seg_3_19_local_g2_7_17379;
  wire seg_3_19_local_g3_2_17382;
  wire seg_3_19_lutff_0_out_13484;
  wire seg_3_19_lutff_1_out_13485;
  wire seg_3_19_lutff_2_out_13486;
  wire seg_3_19_lutff_3_out_13487;
  wire seg_3_19_lutff_4_out_13488;
  wire seg_3_19_lutff_5_out_13489;
  wire seg_3_19_lutff_6_out_13490;
  wire seg_3_19_lutff_7_out_13491;
  wire seg_3_20_glb_netwk_0_5;
  wire seg_3_20_local_g0_2_17481;
  wire seg_3_20_local_g1_6_17493;
  wire seg_3_20_local_g2_0_17495;
  wire seg_3_20_local_g2_5_17500;
  wire seg_3_20_local_g3_1_17504;
  wire seg_3_20_local_g3_3_17506;
  wire seg_3_20_local_g3_4_17507;
  wire seg_3_20_local_g3_7_17510;
  wire seg_3_20_lutff_0_out_13607;
  wire seg_3_20_lutff_1_out_13608;
  wire seg_3_20_lutff_2_out_13609;
  wire seg_3_20_lutff_3_out_13610;
  wire seg_3_20_lutff_4_out_13611;
  wire seg_3_20_lutff_5_out_13612;
  wire seg_3_20_lutff_6_out_13613;
  wire seg_3_20_lutff_7_out_13614;
  wire seg_3_4_sp4_h_r_10_15607;
  wire seg_3_5_sp4_v_t_39_12035;
  wire seg_3_7_glb_netwk_0_5;
  wire seg_3_7_local_g0_7_15887;
  wire seg_3_7_local_g1_5_15893;
  wire seg_3_7_local_g1_7_15895;
  wire seg_3_7_lutff_7_out_12015;
  wire seg_3_7_sp4_v_b_13_11910;
  wire seg_3_7_sp4_v_b_23_11920;
  wire seg_3_7_sp4_v_b_30_12039;
  wire seg_3_8_glb_netwk_0_5;
  wire seg_3_8_local_g1_3_16014;
  wire seg_3_8_local_g1_4_16015;
  wire seg_3_8_local_g1_5_16016;
  wire seg_3_8_lutff_4_out_12135;
  wire seg_3_8_sp4_h_l_46_1816;
  wire seg_3_8_sp4_h_r_7_16106;
  wire seg_3_8_sp4_v_b_19_12039;
  wire seg_3_8_sp4_v_b_5_11913;
  wire seg_4_10_sp4_h_r_1_20175;
  wire seg_4_12_glb_netwk_0_5;
  wire seg_4_12_local_g1_7_20341;
  wire seg_4_12_local_g3_2_20352;
  wire seg_4_12_lutff_2_out_16456;
  wire seg_4_12_sp4_h_r_15_16593;
  wire seg_4_12_sp4_h_r_4_20426;
  wire seg_4_13_glb_netwk_0_5;
  wire seg_4_13_local_g1_4_20461;
  wire seg_4_13_local_g1_5_20462;
  wire seg_4_13_local_g3_5_20478;
  wire seg_4_13_lutff_5_out_16582;
  wire seg_4_13_sp4_h_l_46_2864;
  wire seg_4_13_sp4_v_b_10_16366;
  wire seg_4_13_sp4_v_b_12_16478;
  wire seg_4_13_sp4_v_b_5_16359;
  wire seg_4_14_sp4_h_r_6_20674;
  wire seg_4_17_glb_netwk_0_5;
  wire seg_4_17_local_g0_1_20942;
  wire seg_4_17_local_g3_3_20968;
  wire seg_4_17_lutff_1_out_17070;
  wire seg_4_17_sp4_v_b_27_17095;
  wire seg_4_18_glb_netwk_0_5;
  wire seg_4_18_local_g0_1_21065;
  wire seg_4_18_local_g0_2_21066;
  wire seg_4_18_local_g0_5_21069;
  wire seg_4_18_local_g0_6_21070;
  wire seg_4_18_local_g1_0_21072;
  wire seg_4_18_local_g1_1_21073;
  wire seg_4_18_local_g1_3_21075;
  wire seg_4_18_local_g1_4_21076;
  wire seg_4_18_local_g1_6_21078;
  wire seg_4_18_local_g2_6_21086;
  wire seg_4_18_local_g2_7_21087;
  wire seg_4_18_local_g3_1_21089;
  wire seg_4_18_lutff_0_out_17192;
  wire seg_4_18_lutff_6_out_17198;
  wire seg_4_18_lutff_7_out_17199;
  wire seg_4_18_neigh_op_bot_1_17070;
  wire seg_4_18_neigh_op_lft_2_13363;
  wire seg_4_18_neigh_op_lft_3_13364;
  wire seg_4_18_neigh_op_lft_4_13365;
  wire seg_4_18_neigh_op_lft_5_13366;
  wire seg_4_18_neigh_op_lft_6_13367;
  wire seg_4_18_neigh_op_tnl_1_13485;
  wire seg_4_18_neigh_op_top_1_17316;
  wire seg_4_18_sp4_h_r_4_21164;
  wire seg_4_18_sp4_r_v_b_21_20933;
  wire seg_4_18_sp4_r_v_b_37_21171;
  wire seg_4_18_sp4_r_v_b_5_20805;
  wire seg_4_18_sp4_v_b_14_17095;
  wire seg_4_18_sp4_v_b_6_16977;
  wire seg_4_19_local_g0_2_21189;
  wire seg_4_19_local_g0_3_21190;
  wire seg_4_19_local_g1_0_21195;
  wire seg_4_19_local_g1_1_21196;
  wire seg_4_19_local_g1_2_21197;
  wire seg_4_19_local_g1_4_21199;
  wire seg_4_19_local_g1_7_21202;
  wire seg_4_19_local_g2_0_21203;
  wire seg_4_19_local_g2_7_21210;
  wire seg_4_19_local_g3_0_21211;
  wire seg_4_19_local_g3_5_21216;
  wire seg_4_19_local_g3_7_21218;
  wire seg_4_19_lutff_1_out_17316;
  wire seg_4_19_lutff_2_out_17317;
  wire seg_4_19_lutff_4_out_17319;
  wire seg_4_19_neigh_op_bnl_7_13368;
  wire seg_4_19_neigh_op_lft_0_13484;
  wire seg_4_19_neigh_op_lft_2_13486;
  wire seg_4_19_neigh_op_lft_3_13487;
  wire seg_4_19_neigh_op_lft_7_13491;
  wire seg_4_19_neigh_op_tnl_0_13607;
  wire seg_4_19_neigh_op_tnl_5_13612;
  wire seg_4_19_neigh_op_tnl_7_13614;
  wire seg_4_19_neigh_op_top_1_17439;
  wire seg_4_19_sp4_h_r_24_13619;
  wire seg_4_20_local_g0_3_21313;
  wire seg_4_20_local_g0_6_21316;
  wire seg_4_20_local_g1_1_21319;
  wire seg_4_20_local_g1_4_21322;
  wire seg_4_20_lutff_1_out_17439;
  wire seg_4_20_neigh_op_lft_1_13608;
  wire seg_4_20_neigh_op_lft_3_13610;
  wire seg_4_20_neigh_op_lft_4_13611;
  wire seg_4_20_neigh_op_lft_6_13613;
  wire seg_5_0_span4_vert_13_19048;
  wire seg_5_10_sp4_v_t_40_20313;
  wire seg_5_12_glb_netwk_0_5;
  wire seg_5_12_local_g0_2_24159;
  wire seg_5_12_local_g2_2_24175;
  wire seg_5_12_lutff_2_out_20287;
  wire seg_5_12_neigh_op_lft_2_16456;
  wire seg_5_12_sp4_h_r_4_24257;
  wire seg_5_14_sp4_v_t_40_20805;
  wire seg_5_17_sp4_v_t_37_21171;
  wire seg_5_19_sp4_v_b_8_20933;
  wire seg_5_20_glb_netwk_0_5;
  wire seg_5_20_glb_netwk_3_8;
  wire seg_5_20_local_g1_3_25152;
  wire seg_5_20_sp12_h_r_3_21400;
  wire seg_5_20_sp4_h_r_4_25241;
  wire seg_5_2_sp4_v_t_44_19333;
  wire seg_5_5_glb_netwk_0_5;
  wire seg_5_5_local_g3_7_23327;
  wire seg_5_5_sp4_h_r_0_23390;
  wire seg_5_5_sp4_h_r_31_15737;
  wire seg_5_5_sp4_r_v_b_17_23161;
  wire seg_5_6_sp4_v_t_36_19817;
  wire seg_6_0_glb_netwk_0_5;
  wire seg_6_0_local_g0_2_26539;
  wire seg_6_0_local_g1_2_26547;
  wire seg_6_0_local_g1_6_26551;
  wire seg_6_0_local_g1_6_26551_i1;
  wire seg_6_0_local_g1_6_26551_i2;
  wire seg_6_0_local_g1_6_26551_i3;
  wire seg_6_0_span12_vert_18_26571;
  wire seg_6_0_span4_horz_r_6_22756;
  wire seg_6_0_span4_vert_18_22884;
  wire seg_6_0_span4_vert_32_22900;
  wire seg_6_0_span4_vert_42_22911;
  wire seg_6_10_sp12_v_b_1_26571;
  wire seg_6_13_sp4_h_l_38_12886;
  wire seg_6_17_sp4_v_b_3_24511;
  wire seg_6_28_sp4_h_r_2_29465;
  wire seg_6_2_sp4_h_r_2_26813;
  wire seg_6_2_sp4_v_t_41_23161;
  wire seg_6_31_local_g0_7_29714;
  wire seg_6_31_local_g0_7_29714_i1;
  wire seg_6_31_local_g0_7_29714_i2;
  wire seg_6_31_local_g0_7_29714_i3;
  wire seg_6_31_span4_vert_15_26357;
  wire seg_6_3_sp4_v_b_8_22900;
  wire seg_6_4_sp4_h_l_36_11775;
  wire seg_6_4_sp4_h_r_10_27015;
  wire seg_7_0_glb_netwk_0_5;
  wire seg_7_0_local_g0_6_29743;
  wire seg_7_0_local_g1_2_29747;
  wire seg_7_0_span4_horz_r_14_18925;
  wire seg_7_0_span4_vert_16_26691;
  wire seg_7_0_span4_vert_42_26720;
  wire seg_7_10_sp4_h_r_3_31041;
  wire seg_7_10_sp4_v_b_3_27333;
  wire seg_7_12_glb_netwk_0_5;
  wire seg_7_12_local_g2_3_31207;
  wire seg_7_12_local_g2_4_31208;
  wire seg_7_12_local_g3_1_31213;
  wire seg_7_12_local_g3_2_31214;
  wire seg_7_12_lutff_2_out_27687;
  wire seg_7_12_lutff_3_out_27688;
  wire seg_7_12_sp4_h_r_10_31284;
  wire seg_7_12_sp4_h_r_28_24257;
  wire seg_7_12_sp4_h_r_41_20426;
  wire seg_7_12_sp4_v_b_9_27543;
  wire seg_7_1_local_g2_3_29814;
  wire seg_7_1_local_g3_7_29826;
  wire seg_7_1_neigh_op_tnr_3_29884;
  wire seg_7_1_neigh_op_tnr_7_29888;
  wire seg_7_28_sp12_h_r_6_22385;
  wire seg_7_2_sp4_v_b_5_26691;
  wire seg_7_4_sp4_h_r_7_30307;
  wire seg_7_8_sp4_v_b_1_27127;
  wire seg_8_0_span4_vert_37_29936;
  wire seg_8_10_glb_netwk_0_5;
  wire seg_8_10_local_g0_2_34775;
  wire seg_8_10_local_g0_4_34777;
  wire seg_8_10_local_g0_5_34778;
  wire seg_8_10_local_g0_6_34779;
  wire seg_8_10_local_g1_5_34786;
  wire seg_8_10_local_g3_2_34799;
  wire seg_8_10_local_g3_3_34800;
  wire seg_8_10_local_g3_4_34801;
  wire seg_8_10_lutff_2_out_30903;
  wire seg_8_10_lutff_3_out_30904;
  wire seg_8_10_lutff_4_out_30905;
  wire seg_8_10_lutff_5_out_30906;
  wire seg_8_10_lutff_6_out_30907;
  wire seg_8_10_neigh_op_top_5_31029;
  wire seg_8_10_sp12_v_b_14_34250;
  wire seg_8_10_sp4_h_r_14_31041;
  wire seg_8_10_sp4_h_r_20_31047;
  wire seg_8_10_sp4_h_r_30_27633;
  wire seg_8_10_sp4_h_r_46_24008;
  wire seg_8_10_sp4_v_b_1_30679;
  wire seg_8_10_sp4_v_b_26_30928;
  wire seg_8_11_glb_netwk_0_5;
  wire seg_8_11_local_g0_2_34898;
  wire seg_8_11_local_g0_5_34901;
  wire seg_8_11_local_g3_5_34925;
  wire seg_8_11_lutff_5_out_31029;
  wire seg_8_11_sp12_v_b_13_34250;
  wire seg_8_11_sp4_v_b_18_30931;
  wire seg_8_12_glb_netwk_0_5;
  wire seg_8_12_local_g0_1_35020;
  wire seg_8_12_local_g0_4_35023;
  wire seg_8_12_local_g3_2_35045;
  wire seg_8_12_lutff_1_out_31148;
  wire seg_8_12_sp12_v_b_2_33722;
  wire seg_8_12_sp4_h_r_2_35117;
  wire seg_8_12_sp4_r_v_b_28_35007;
  wire seg_8_12_sp4_v_b_2_30928;
  wire seg_8_13_sp12_v_b_1_33722;
  wire seg_8_14_sp4_v_b_1_31171;
  wire seg_8_17_glb_netwk_0_5;
  wire seg_8_17_local_g2_1_35651;
  wire seg_8_17_sp4_h_r_26_28343;
  wire seg_8_17_sp4_h_r_33_28350;
  wire seg_8_17_sp4_r_v_b_43_35747;
  wire seg_8_18_sp4_h_l_41_21164;
  wire seg_8_23_glb_netwk_0_5;
  wire seg_8_23_local_g0_4_36376;
  wire seg_8_23_local_g2_5_36393;
  wire seg_8_23_local_g3_5_36401;
  wire seg_8_23_lutff_5_out_32505;
  wire seg_8_23_sp12_v_b_5_35234;
  wire seg_8_23_sp4_h_r_4_36472;
  wire seg_8_23_sp4_v_b_26_32527;
  wire seg_8_23_sp4_v_t_41_32775;
  wire seg_8_24_glb_netwk_0_5;
  wire seg_8_24_local_g0_2_36497;
  wire seg_8_24_local_g1_5_36508;
  wire seg_8_24_local_g2_6_36517;
  wire seg_8_24_lutff_6_out_32629;
  wire seg_8_24_sp4_v_b_18_32530;
  wire seg_8_24_sp4_v_b_3_32403;
  wire seg_8_24_sp4_v_b_5_32405;
  wire seg_8_24_sp4_v_t_44_32901;
  wire seg_8_25_glb_netwk_0_5;
  wire seg_8_25_local_g0_3_36621;
  wire seg_8_25_local_g0_4_36622;
  wire seg_8_25_local_g0_6_36624;
  wire seg_8_25_local_g1_2_36628;
  wire seg_8_25_local_g1_4_36630;
  wire seg_8_25_local_g1_7_36633;
  wire seg_8_25_local_g2_2_36636;
  wire seg_8_25_local_g3_5_36647;
  wire seg_8_25_lutff_2_out_32748;
  wire seg_8_25_lutff_3_out_32749;
  wire seg_8_25_lutff_4_out_32750;
  wire seg_8_25_lutff_5_out_32751;
  wire seg_8_25_lutff_7_out_32753;
  wire seg_8_25_neigh_op_bot_6_32629;
  wire seg_8_25_sp12_v_b_1_35234;
  wire seg_8_25_sp4_h_r_12_32882;
  wire seg_8_25_sp4_h_r_2_36716;
  wire seg_8_25_sp4_r_v_b_29_36605;
  wire seg_8_25_sp4_v_b_28_32775;
  wire seg_8_25_sp4_v_b_2_32527;
  wire seg_8_25_sp4_v_b_44_32901;
  wire seg_8_28_sp4_v_b_11_32903;
  wire seg_8_2_glb_netwk_0_5;
  wire seg_8_2_local_g0_2_33791;
  wire seg_8_2_local_g1_0_33797;
  wire seg_8_2_local_g1_5_33802;
  wire seg_8_2_local_g1_6_33803;
  wire seg_8_2_local_g2_0_33805;
  wire seg_8_2_local_g3_1_33814;
  wire seg_8_2_local_g3_2_33815;
  wire seg_8_2_local_g3_3_33816;
  wire seg_8_2_local_g3_4_33817;
  wire seg_8_2_lutff_1_out_29882;
  wire seg_8_2_lutff_2_out_29883;
  wire seg_8_2_lutff_3_out_29884;
  wire seg_8_2_lutff_6_out_29887;
  wire seg_8_2_lutff_7_out_29888;
  wire seg_8_2_neigh_op_rgt_0_33712;
  wire seg_8_2_neigh_op_tnr_1_33872;
  wire seg_8_2_neigh_op_tnr_2_33873;
  wire seg_8_2_neigh_op_tnr_4_33875;
  wire seg_8_2_neigh_op_top_5_30045;
  wire seg_8_2_sp4_h_r_16_30059;
  wire seg_8_2_sp4_h_r_26_26813;
  wire seg_8_2_sp4_r_v_b_43_33902;
  wire seg_8_2_sp4_v_b_24_29936;
  wire seg_8_30_sp4_v_t_36_37347;
  wire seg_8_31_glb_netwk_0_5;
  wire seg_8_31_io_1_D_IN_0_33486;
  wire seg_8_31_local_g0_7_37376;
  wire seg_8_31_local_g1_5_37382;
  wire seg_8_31_logic_op_bnr_7_37199;
  wire seg_8_31_span12_vert_13_36710;
  wire seg_8_31_span4_horz_r_6_33556;
  wire seg_8_31_span4_vert_36_37347;
  wire seg_8_3_glb_netwk_0_5;
  wire seg_8_3_local_g0_0_33912;
  wire seg_8_3_local_g0_2_33914;
  wire seg_8_3_local_g0_4_33916;
  wire seg_8_3_local_g1_6_33926;
  wire seg_8_3_local_g2_1_33929;
  wire seg_8_3_local_g2_4_33932;
  wire seg_8_3_local_g3_2_33938;
  wire seg_8_3_local_g3_5_33941;
  wire seg_8_3_lutff_4_out_30044;
  wire seg_8_3_lutff_5_out_30045;
  wire seg_8_3_lutff_6_out_30046;
  wire seg_8_3_neigh_op_rgt_1_33872;
  wire seg_8_3_neigh_op_rgt_2_33873;
  wire seg_8_3_neigh_op_rgt_4_33875;
  wire seg_8_3_sp4_h_r_18_30184;
  wire seg_8_3_sp4_h_r_30_26919;
  wire seg_8_3_sp4_r_v_b_19_33774;
  wire seg_8_3_sp4_r_v_b_24_33896;
  wire seg_8_4_lutff_1_out_30164;
  wire seg_8_4_sp12_v_b_18_33722;
  wire seg_8_4_sp4_h_r_18_30307;
  wire seg_8_4_sp4_h_r_2_34133;
  wire seg_8_4_sp4_h_r_34_27015;
  wire seg_8_4_sp4_r_v_b_35_34028;
  wire seg_8_4_sp4_r_v_b_3_33768;
  wire seg_8_4_sp4_v_b_34_30198;
  wire seg_8_6_sp4_v_b_10_30198;
  wire seg_9_10_glb_netwk_0_5;
  wire seg_9_10_local_g0_6_38610;
  wire seg_9_10_local_g2_2_38622;
  wire seg_9_10_local_g2_7_38627;
  wire seg_9_10_local_g3_2_38630;
  wire seg_9_10_local_g3_4_38632;
  wire seg_9_10_local_g3_7_38635;
  wire seg_9_10_lutff_1_out_34733;
  wire seg_9_10_lutff_2_out_34734;
  wire seg_9_10_lutff_4_out_34736;
  wire seg_9_10_lutff_7_out_34739;
  wire seg_9_10_sp12_h_r_6_27622;
  wire seg_9_10_sp4_h_l_40_24012;
  wire seg_9_10_sp4_h_l_46_24008;
  wire seg_9_10_sp4_h_r_12_34868;
  wire seg_9_10_sp4_h_r_2_38702;
  wire seg_9_10_sp4_r_v_b_10_38352;
  wire seg_9_10_sp4_r_v_b_23_38475;
  wire seg_9_10_sp4_r_v_b_41_38715;
  wire seg_9_11_glb_netwk_0_5;
  wire seg_9_11_glb_netwk_1_6;
  wire seg_9_11_local_g2_2_38745;
  wire seg_9_11_lutff_5_out_34860;
  wire seg_9_11_sp4_h_r_10_38823;
  wire seg_9_11_sp4_r_v_b_10_38475;
  wire seg_9_12_glb_netwk_0_5;
  wire seg_9_12_local_g1_6_38864;
  wire seg_9_12_local_g2_2_38868;
  wire seg_9_12_sp4_h_r_34_31284;
  wire seg_9_12_sp4_r_v_b_35_38843;
  wire seg_9_12_sp4_r_v_b_3_38589;
  wire seg_9_12_sp4_v_b_2_34759;
  wire seg_9_12_sp4_v_b_6_34763;
  wire seg_9_17_sp4_h_l_40_24873;
  wire seg_9_18_glb_netwk_0_5;
  wire seg_9_18_glb_netwk_1_6;
  wire seg_9_18_local_g2_5_39609;
  wire seg_9_18_local_g2_6_39610;
  wire seg_9_18_neigh_op_tnr_5_39675;
  wire seg_9_18_neigh_op_tnr_6_39676;
  wire seg_9_18_sp4_h_r_2_39686;
  wire seg_9_18_sp4_r_v_b_11_39335;
  wire seg_9_19_sp4_h_l_45_25122;
  wire seg_9_20_sp4_h_l_41_25241;
  wire seg_9_20_sp4_v_b_6_35747;
  wire seg_9_23_sp4_v_t_40_36605;
  wire seg_9_24_sp4_v_b_2_36235;
  wire seg_9_27_glb_netwk_0_5;
  wire seg_9_27_local_g0_1_40696;
  wire seg_9_27_local_g1_3_40706;
  wire seg_9_27_local_g2_4_40715;
  wire seg_9_27_local_g2_7_40718;
  wire seg_9_27_local_g3_0_40719;
  wire seg_9_27_local_g3_2_40721;
  wire seg_9_27_lutff_1_out_36824;
  wire seg_9_27_lutff_5_out_36828;
  wire seg_9_27_lutff_7_out_36830;
  wire seg_9_27_neigh_op_rgt_2_40656;
  wire seg_9_27_sp4_r_v_b_16_40559;
  wire seg_9_27_sp4_r_v_b_27_40680;
  wire seg_9_27_sp4_r_v_b_36_40801;
  wire seg_9_28_glb_netwk_0_5;
  wire seg_9_28_local_g0_0_40818;
  wire seg_9_28_local_g0_2_40820;
  wire seg_9_28_local_g0_5_40823;
  wire seg_9_28_local_g0_7_40825;
  wire seg_9_28_local_g1_0_40826;
  wire seg_9_28_local_g1_2_40828;
  wire seg_9_28_local_g1_5_40831;
  wire seg_9_28_local_g1_7_40833;
  wire seg_9_28_local_g2_2_40836;
  wire seg_9_28_local_g2_3_40837;
  wire seg_9_28_local_g2_5_40839;
  wire seg_9_28_lutff_2_out_36948;
  wire seg_9_28_lutff_5_out_36951;
  wire seg_9_28_neigh_op_bnr_7_40661;
  wire seg_9_28_neigh_op_bot_5_36828;
  wire seg_9_28_neigh_op_bot_7_36830;
  wire seg_9_28_neigh_op_rgt_3_40780;
  wire seg_9_28_neigh_op_top_5_37074;
  wire seg_9_28_sp4_h_r_16_37088;
  wire seg_9_28_sp4_h_r_34_33252;
  wire seg_9_28_sp4_v_b_2_36727;
  wire seg_9_28_sp4_v_b_44_37101;
  wire seg_9_29_local_g0_0_40941;
  wire seg_9_29_local_g1_1_40950;
  wire seg_9_29_local_g2_0_40957;
  wire seg_9_29_local_g2_3_40960;
  wire seg_9_29_local_g2_4_40961;
  wire seg_9_29_local_g2_5_40962;
  wire seg_9_29_local_g3_0_40965;
  wire seg_9_29_local_g3_5_40970;
  wire seg_9_29_lutff_0_out_37069;
  wire seg_9_29_lutff_3_out_37072;
  wire seg_9_29_lutff_5_out_37074;
  wire seg_9_29_neigh_op_rgt_0_40900;
  wire seg_9_29_neigh_op_rgt_5_40905;
  wire seg_9_29_neigh_op_tnr_3_41026;
  wire seg_9_29_neigh_op_tnr_4_41027;
  wire seg_9_29_sp4_h_r_38_29568;
  wire seg_9_29_sp4_r_v_b_1_40678;
  wire seg_9_2_glb_netwk_0_5;
  wire seg_9_2_local_g0_1_37621;
  wire seg_9_2_local_g0_2_37622;
  wire seg_9_2_local_g0_3_37623;
  wire seg_9_2_local_g0_4_37624;
  wire seg_9_2_local_g0_7_37627;
  wire seg_9_2_local_g1_3_37631;
  wire seg_9_2_local_g1_4_37632;
  wire seg_9_2_local_g1_5_37633;
  wire seg_9_2_local_g1_7_37635;
  wire seg_9_2_local_g2_1_37637;
  wire seg_9_2_local_g2_2_37638;
  wire seg_9_2_local_g2_3_37639;
  wire seg_9_2_local_g2_4_37640;
  wire seg_9_2_local_g2_6_37642;
  wire seg_9_2_local_g2_7_37643;
  wire seg_9_2_local_g3_2_37646;
  wire seg_9_2_local_g3_3_37647;
  wire seg_9_2_local_g3_4_37648;
  wire seg_9_2_local_g3_5_37649;
  wire seg_9_2_local_g3_6_37650;
  wire seg_9_2_local_g3_7_37651;
  wire seg_9_2_lutff_0_out_33712;
  wire seg_9_2_lutff_1_out_33713;
  wire seg_9_2_lutff_2_out_33714;
  wire seg_9_2_lutff_3_out_33715;
  wire seg_9_2_lutff_4_out_33716;
  wire seg_9_2_lutff_5_out_33717;
  wire seg_9_2_lutff_6_out_33718;
  wire seg_9_2_lutff_7_out_33719;
  wire seg_9_2_neigh_op_lft_3_29884;
  wire seg_9_2_neigh_op_rgt_6_37549;
  wire seg_9_2_neigh_op_rgt_7_37550;
  wire seg_9_2_neigh_op_tnl_5_30045;
  wire seg_9_2_neigh_op_tnr_2_37704;
  wire seg_9_2_neigh_op_tnr_3_37705;
  wire seg_9_2_neigh_op_tnr_4_37706;
  wire seg_9_2_neigh_op_tnr_6_37708;
  wire seg_9_2_neigh_op_top_1_33872;
  wire seg_9_2_neigh_op_top_2_33873;
  wire seg_9_2_neigh_op_top_4_33875;
  wire seg_9_2_neigh_op_top_7_33878;
  wire seg_9_2_sp4_h_r_44_26820;
  wire seg_9_2_sp4_v_b_27_33768;
  wire seg_9_2_sp4_v_t_46_34028;
  wire seg_9_30_glb_netwk_0_5;
  wire seg_9_30_local_g0_0_41064;
  wire seg_9_30_local_g0_4_41068;
  wire seg_9_30_local_g1_0_41072;
  wire seg_9_30_local_g1_5_41077;
  wire seg_9_30_local_g2_2_41082;
  wire seg_9_30_local_g2_3_41083;
  wire seg_9_30_local_g2_4_41084;
  wire seg_9_30_local_g3_6_41094;
  wire seg_9_30_lutff_0_out_37192;
  wire seg_9_30_lutff_5_out_37197;
  wire seg_9_30_lutff_7_out_37199;
  wire seg_9_30_neigh_op_bnr_0_40900;
  wire seg_9_30_neigh_op_bnr_5_40905;
  wire seg_9_30_neigh_op_rgt_3_41026;
  wire seg_9_30_neigh_op_rgt_4_41027;
  wire seg_9_30_neigh_op_tnl_6_33486;
  wire seg_9_30_sp4_v_b_20_37101;
  wire seg_9_30_sp4_v_b_26_37219;
  wire seg_9_3_glb_netwk_0_5;
  wire seg_9_3_local_g0_5_37748;
  wire seg_9_3_local_g0_6_37749;
  wire seg_9_3_local_g1_1_37752;
  wire seg_9_3_local_g1_3_37754;
  wire seg_9_3_local_g1_4_37755;
  wire seg_9_3_local_g1_5_37756;
  wire seg_9_3_local_g1_6_37757;
  wire seg_9_3_local_g2_0_37759;
  wire seg_9_3_local_g2_1_37760;
  wire seg_9_3_local_g2_4_37763;
  wire seg_9_3_local_g2_5_37764;
  wire seg_9_3_local_g2_7_37766;
  wire seg_9_3_local_g3_1_37768;
  wire seg_9_3_local_g3_2_37769;
  wire seg_9_3_local_g3_3_37770;
  wire seg_9_3_lutff_0_out_33871;
  wire seg_9_3_lutff_1_out_33872;
  wire seg_9_3_lutff_2_out_33873;
  wire seg_9_3_lutff_3_out_33874;
  wire seg_9_3_lutff_4_out_33875;
  wire seg_9_3_lutff_5_out_33876;
  wire seg_9_3_lutff_6_out_33877;
  wire seg_9_3_lutff_7_out_33878;
  wire seg_9_3_neigh_op_bnl_1_29882;
  wire seg_9_3_neigh_op_bot_6_33718;
  wire seg_9_3_neigh_op_lft_5_30045;
  wire seg_9_3_neigh_op_top_5_33999;
  wire seg_9_3_sp4_v_b_19_33774;
  wire seg_9_3_sp4_v_b_24_33896;
  wire seg_9_4_glb_netwk_0_5;
  wire seg_9_4_local_g0_0_37866;
  wire seg_9_4_local_g0_3_37869;
  wire seg_9_4_local_g1_3_37877;
  wire seg_9_4_local_g2_1_37883;
  wire seg_9_4_local_g3_5_37895;
  wire seg_9_4_lutff_1_out_33995;
  wire seg_9_4_lutff_5_out_33999;
  wire seg_9_4_neigh_op_bnl_5_30045;
  wire seg_9_4_neigh_op_bot_0_33871;
  wire seg_9_4_sp4_h_r_3_37965;
  wire seg_9_4_sp4_v_b_16_33899;
  wire seg_9_4_sp4_v_b_19_33902;
  wire seg_9_4_sp4_v_b_3_33768;
  wire seg_9_4_sp4_v_t_47_34275;
  wire seg_9_5_glb_netwk_0_5;
  wire seg_9_5_local_g1_3_38000;
  wire seg_9_5_local_g3_1_38014;
  wire seg_9_5_neigh_op_bnl_1_30164;
  wire seg_9_5_sp4_h_l_37_23390;
  wire seg_9_5_sp4_h_r_11_38086;
  wire seg_9_5_sp4_r_v_b_23_37860;
  wire seg_9_5_sp4_v_b_5_33899;
  wire seg_9_6_sp4_v_b_11_34028;
  wire seg_9_8_local_g0_6_38364;
  wire seg_9_8_local_g1_1_38367;
  wire seg_9_8_local_g1_7_38373;
  wire seg_9_8_local_g2_2_38376;
  wire seg_9_8_local_g2_6_38380;
  wire seg_9_8_local_g3_0_38382;
  wire seg_9_8_local_g3_1_38383;
  wire seg_9_8_local_g3_4_38386;
  wire seg_9_8_lutff_5_out_34491;
  wire seg_9_8_lutff_6_out_34492;
  wire seg_9_8_lutff_7_out_34493;
  wire seg_9_8_neigh_op_rgt_2_38319;
  wire seg_9_8_neigh_op_rgt_4_38321;
  wire seg_9_8_neigh_op_rgt_6_38323;
  wire seg_9_8_sp4_h_r_15_34625;
  wire seg_9_8_sp4_h_r_17_34627;
  wire seg_9_8_sp4_h_r_24_30790;
  wire seg_9_8_sp4_r_v_b_16_38222;
  wire seg_9_8_sp4_r_v_b_17_38223;
  wire seg_9_8_sp4_r_v_b_21_38227;
  wire seg_9_8_sp4_r_v_b_23_38229;
  wire seg_9_8_sp4_v_b_14_34389;
  wire seg_9_8_sp4_v_b_6_34271;
  wire seg_9_8_sp4_v_t_39_34759;
  wire seg_9_9_sp4_h_r_10_38577;
  wire t0;
  wire t10;
  wire t109;
  wire t11;
  wire t113;
  wire t115;
  wire t120;
  wire t122;
  wire t13;
  wire t138;
  wire t140;
  wire t2;
  wire t219;
  wire t245;
  wire t247;
  wire t251;
  wire t253;
  wire t254;
  wire t256;
  wire t285;
  wire t315;
  wire t317;
  wire t399;
  wire t450;
  wire t452;
  wire t455;
  wire t458;
  wire t46;
  wire t48;
  wire t50;
  wire t52;
  wire t55;
  wire t57;
  wire t630;
  wire t67;
  wire t69;
  wire t735;
  wire t753;
  wire t755;
  wire t8;
  wire t81;
  wire t83;
  assign net_10 = seg_22_16_glb_netwk_5_10;
  assign net_11 = seg_22_16_glb_netwk_6_11;
  assign net_12178 = seg_2_8_local_g0_6_12178;
  assign net_12179 = seg_2_8_local_g0_7_12179;
  assign net_12185 = seg_2_8_local_g1_5_12185;
  assign net_12191 = seg_2_8_local_g2_3_12191;
  assign net_12192 = seg_2_8_local_g2_4_12192;
  assign net_12198 = seg_2_8_local_g3_2_12198;
  assign net_12200 = seg_2_8_local_g3_4_12200;
  assign net_12201 = seg_2_8_local_g3_5_12201;
  assign net_13545 = seg_2_19_local_g2_4_13545;
  assign net_13551 = seg_2_19_local_g3_2_13551;
  assign net_13554 = seg_2_19_local_g3_5_13554;
  assign net_13555 = seg_2_19_local_g3_6_13555;
  assign net_15887 = seg_3_7_local_g0_7_15887;
  assign net_15893 = seg_3_7_local_g1_5_15893;
  assign net_15895 = seg_3_7_local_g1_7_15895;
  assign net_16014 = seg_3_8_local_g1_3_16014;
  assign net_16015 = seg_3_8_local_g1_4_16015;
  assign net_16016 = seg_3_8_local_g1_5_16016;
  assign net_16620 = seg_3_13_local_g0_2_16620;
  assign net_16628 = seg_3_13_local_g1_2_16628;
  assign net_16631 = seg_3_13_local_g1_5_16631;
  assign net_16632 = seg_3_13_local_g1_6_16632;
  assign net_16639 = seg_3_13_local_g2_5_16639;
  assign net_16645 = seg_3_13_local_g3_3_16645;
  assign net_16646 = seg_3_13_local_g3_4_16646;
  assign net_16647 = seg_3_13_local_g3_5_16647;
  assign net_16759 = seg_3_14_local_g2_2_16759;
  assign net_16768 = seg_3_14_local_g3_3_16768;
  assign net_16770 = seg_3_14_local_g3_5_16770;
  assign net_17237 = seg_3_18_local_g0_4_17237;
  assign net_17238 = seg_3_18_local_g0_5_17238;
  assign net_17239 = seg_3_18_local_g0_6_17239;
  assign net_17242 = seg_3_18_local_g1_1_17242;
  assign net_17251 = seg_3_18_local_g2_2_17251;
  assign net_17252 = seg_3_18_local_g2_3_17252;
  assign net_17256 = seg_3_18_local_g2_7_17256;
  assign net_17264 = seg_3_18_local_g3_7_17264;
  assign net_17357 = seg_3_19_local_g0_1_17357;
  assign net_17362 = seg_3_19_local_g0_6_17362;
  assign net_17364 = seg_3_19_local_g1_0_17364;
  assign net_17367 = seg_3_19_local_g1_3_17367;
  assign net_17376 = seg_3_19_local_g2_4_17376;
  assign net_17377 = seg_3_19_local_g2_5_17377;
  assign net_17379 = seg_3_19_local_g2_7_17379;
  assign net_17382 = seg_3_19_local_g3_2_17382;
  assign net_17481 = seg_3_20_local_g0_2_17481;
  assign net_17493 = seg_3_20_local_g1_6_17493;
  assign net_17495 = seg_3_20_local_g2_0_17495;
  assign net_17500 = seg_3_20_local_g2_5_17500;
  assign net_17504 = seg_3_20_local_g3_1_17504;
  assign net_17506 = seg_3_20_local_g3_3_17506;
  assign net_17507 = seg_3_20_local_g3_4_17507;
  assign net_17510 = seg_3_20_local_g3_7_17510;
  assign net_20341 = seg_4_12_local_g1_7_20341;
  assign net_20352 = seg_4_12_local_g3_2_20352;
  assign net_20461 = seg_4_13_local_g1_4_20461;
  assign net_20462 = seg_4_13_local_g1_5_20462;
  assign net_20478 = seg_4_13_local_g3_5_20478;
  assign net_20942 = seg_4_17_local_g0_1_20942;
  assign net_20968 = seg_4_17_local_g3_3_20968;
  assign net_21065 = seg_4_18_local_g0_1_21065;
  assign net_21066 = seg_4_18_local_g0_2_21066;
  assign net_21069 = seg_4_18_local_g0_5_21069;
  assign net_21070 = seg_4_18_local_g0_6_21070;
  assign net_21072 = seg_4_18_local_g1_0_21072;
  assign net_21073 = seg_4_18_local_g1_1_21073;
  assign net_21075 = seg_4_18_local_g1_3_21075;
  assign net_21076 = seg_4_18_local_g1_4_21076;
  assign net_21078 = seg_4_18_local_g1_6_21078;
  assign net_21086 = seg_4_18_local_g2_6_21086;
  assign net_21087 = seg_4_18_local_g2_7_21087;
  assign net_21089 = seg_4_18_local_g3_1_21089;
  assign net_21189 = seg_4_19_local_g0_2_21189;
  assign net_21190 = seg_4_19_local_g0_3_21190;
  assign net_21195 = seg_4_19_local_g1_0_21195;
  assign net_21196 = seg_4_19_local_g1_1_21196;
  assign net_21197 = seg_4_19_local_g1_2_21197;
  assign net_21199 = seg_4_19_local_g1_4_21199;
  assign net_21202 = seg_4_19_local_g1_7_21202;
  assign net_21203 = seg_4_19_local_g2_0_21203;
  assign net_21210 = seg_4_19_local_g2_7_21210;
  assign net_21211 = seg_4_19_local_g3_0_21211;
  assign net_21216 = seg_4_19_local_g3_5_21216;
  assign net_21218 = seg_4_19_local_g3_7_21218;
  assign net_21313 = seg_4_20_local_g0_3_21313;
  assign net_21316 = seg_4_20_local_g0_6_21316;
  assign net_21319 = seg_4_20_local_g1_1_21319;
  assign net_21322 = seg_4_20_local_g1_4_21322;
  assign net_23327 = seg_5_5_local_g3_7_23327;
  assign net_24159 = seg_5_12_local_g0_2_24159;
  assign net_24175 = seg_5_12_local_g2_2_24175;
  assign net_25152 = seg_5_20_local_g1_3_25152;
  assign net_26539 = seg_6_0_local_g0_2_26539;
  assign net_26547 = seg_6_0_local_g1_2_26547;
  assign net_29743 = seg_7_0_local_g0_6_29743;
  assign net_29747 = seg_7_0_local_g1_2_29747;
  assign net_29814 = seg_7_1_local_g2_3_29814;
  assign net_29826 = seg_7_1_local_g3_7_29826;
  assign net_31207 = seg_7_12_local_g2_3_31207;
  assign net_31208 = seg_7_12_local_g2_4_31208;
  assign net_31213 = seg_7_12_local_g3_1_31213;
  assign net_31214 = seg_7_12_local_g3_2_31214;
  assign net_33791 = seg_8_2_local_g0_2_33791;
  assign net_33797 = seg_8_2_local_g1_0_33797;
  assign net_33802 = seg_8_2_local_g1_5_33802;
  assign net_33803 = seg_8_2_local_g1_6_33803;
  assign net_33805 = seg_8_2_local_g2_0_33805;
  assign net_33814 = seg_8_2_local_g3_1_33814;
  assign net_33815 = seg_8_2_local_g3_2_33815;
  assign net_33816 = seg_8_2_local_g3_3_33816;
  assign net_33817 = seg_8_2_local_g3_4_33817;
  assign net_33912 = seg_8_3_local_g0_0_33912;
  assign net_33914 = seg_8_3_local_g0_2_33914;
  assign net_33916 = seg_8_3_local_g0_4_33916;
  assign net_33926 = seg_8_3_local_g1_6_33926;
  assign net_33929 = seg_8_3_local_g2_1_33929;
  assign net_33932 = seg_8_3_local_g2_4_33932;
  assign net_33938 = seg_8_3_local_g3_2_33938;
  assign net_33941 = seg_8_3_local_g3_5_33941;
  assign net_34775 = seg_8_10_local_g0_2_34775;
  assign net_34777 = seg_8_10_local_g0_4_34777;
  assign net_34778 = seg_8_10_local_g0_5_34778;
  assign net_34779 = seg_8_10_local_g0_6_34779;
  assign net_34786 = seg_8_10_local_g1_5_34786;
  assign net_34799 = seg_8_10_local_g3_2_34799;
  assign net_34800 = seg_8_10_local_g3_3_34800;
  assign net_34801 = seg_8_10_local_g3_4_34801;
  assign net_34898 = seg_8_11_local_g0_2_34898;
  assign net_34901 = seg_8_11_local_g0_5_34901;
  assign net_34925 = seg_8_11_local_g3_5_34925;
  assign net_35020 = seg_8_12_local_g0_1_35020;
  assign net_35023 = seg_8_12_local_g0_4_35023;
  assign net_35045 = seg_8_12_local_g3_2_35045;
  assign net_35651 = seg_8_17_local_g2_1_35651;
  assign net_36376 = seg_8_23_local_g0_4_36376;
  assign net_36393 = seg_8_23_local_g2_5_36393;
  assign net_36401 = seg_8_23_local_g3_5_36401;
  assign net_36497 = seg_8_24_local_g0_2_36497;
  assign net_36508 = seg_8_24_local_g1_5_36508;
  assign net_36517 = seg_8_24_local_g2_6_36517;
  assign net_36621 = seg_8_25_local_g0_3_36621;
  assign net_36622 = seg_8_25_local_g0_4_36622;
  assign net_36624 = seg_8_25_local_g0_6_36624;
  assign net_36628 = seg_8_25_local_g1_2_36628;
  assign net_36630 = seg_8_25_local_g1_4_36630;
  assign net_36633 = seg_8_25_local_g1_7_36633;
  assign net_36636 = seg_8_25_local_g2_2_36636;
  assign net_36647 = seg_8_25_local_g3_5_36647;
  assign net_37376 = seg_8_31_local_g0_7_37376;
  assign net_37382 = seg_8_31_local_g1_5_37382;
  assign net_37621 = seg_9_2_local_g0_1_37621;
  assign net_37622 = seg_9_2_local_g0_2_37622;
  assign net_37623 = seg_9_2_local_g0_3_37623;
  assign net_37624 = seg_9_2_local_g0_4_37624;
  assign net_37627 = seg_9_2_local_g0_7_37627;
  assign net_37631 = seg_9_2_local_g1_3_37631;
  assign net_37632 = seg_9_2_local_g1_4_37632;
  assign net_37633 = seg_9_2_local_g1_5_37633;
  assign net_37635 = seg_9_2_local_g1_7_37635;
  assign net_37637 = seg_9_2_local_g2_1_37637;
  assign net_37638 = seg_9_2_local_g2_2_37638;
  assign net_37639 = seg_9_2_local_g2_3_37639;
  assign net_37640 = seg_9_2_local_g2_4_37640;
  assign net_37642 = seg_9_2_local_g2_6_37642;
  assign net_37643 = seg_9_2_local_g2_7_37643;
  assign net_37646 = seg_9_2_local_g3_2_37646;
  assign net_37647 = seg_9_2_local_g3_3_37647;
  assign net_37648 = seg_9_2_local_g3_4_37648;
  assign net_37649 = seg_9_2_local_g3_5_37649;
  assign net_37650 = seg_9_2_local_g3_6_37650;
  assign net_37651 = seg_9_2_local_g3_7_37651;
  assign net_37748 = seg_9_3_local_g0_5_37748;
  assign net_37749 = seg_9_3_local_g0_6_37749;
  assign net_37752 = seg_9_3_local_g1_1_37752;
  assign net_37754 = seg_9_3_local_g1_3_37754;
  assign net_37755 = seg_9_3_local_g1_4_37755;
  assign net_37756 = seg_9_3_local_g1_5_37756;
  assign net_37757 = seg_9_3_local_g1_6_37757;
  assign net_37759 = seg_9_3_local_g2_0_37759;
  assign net_37760 = seg_9_3_local_g2_1_37760;
  assign net_37763 = seg_9_3_local_g2_4_37763;
  assign net_37764 = seg_9_3_local_g2_5_37764;
  assign net_37766 = seg_9_3_local_g2_7_37766;
  assign net_37768 = seg_9_3_local_g3_1_37768;
  assign net_37769 = seg_9_3_local_g3_2_37769;
  assign net_37770 = seg_9_3_local_g3_3_37770;
  assign net_37866 = seg_9_4_local_g0_0_37866;
  assign net_37869 = seg_9_4_local_g0_3_37869;
  assign net_37877 = seg_9_4_local_g1_3_37877;
  assign net_37883 = seg_9_4_local_g2_1_37883;
  assign net_37895 = seg_9_4_local_g3_5_37895;
  assign net_38000 = seg_9_5_local_g1_3_38000;
  assign net_38014 = seg_9_5_local_g3_1_38014;
  assign net_38364 = seg_9_8_local_g0_6_38364;
  assign net_38367 = seg_9_8_local_g1_1_38367;
  assign net_38373 = seg_9_8_local_g1_7_38373;
  assign net_38376 = seg_9_8_local_g2_2_38376;
  assign net_38380 = seg_9_8_local_g2_6_38380;
  assign net_38382 = seg_9_8_local_g3_0_38382;
  assign net_38383 = seg_9_8_local_g3_1_38383;
  assign net_38386 = seg_9_8_local_g3_4_38386;
  assign net_38610 = seg_9_10_local_g0_6_38610;
  assign net_38622 = seg_9_10_local_g2_2_38622;
  assign net_38627 = seg_9_10_local_g2_7_38627;
  assign net_38630 = seg_9_10_local_g3_2_38630;
  assign net_38632 = seg_9_10_local_g3_4_38632;
  assign net_38635 = seg_9_10_local_g3_7_38635;
  assign net_38745 = seg_9_11_local_g2_2_38745;
  assign net_38864 = seg_9_12_local_g1_6_38864;
  assign net_38868 = seg_9_12_local_g2_2_38868;
  assign net_39609 = seg_9_18_local_g2_5_39609;
  assign net_39610 = seg_9_18_local_g2_6_39610;
  assign net_40696 = seg_9_27_local_g0_1_40696;
  assign net_40706 = seg_9_27_local_g1_3_40706;
  assign net_40715 = seg_9_27_local_g2_4_40715;
  assign net_40718 = seg_9_27_local_g2_7_40718;
  assign net_40719 = seg_9_27_local_g3_0_40719;
  assign net_40721 = seg_9_27_local_g3_2_40721;
  assign net_40818 = seg_9_28_local_g0_0_40818;
  assign net_40820 = seg_9_28_local_g0_2_40820;
  assign net_40823 = seg_9_28_local_g0_5_40823;
  assign net_40825 = seg_9_28_local_g0_7_40825;
  assign net_40826 = seg_9_28_local_g1_0_40826;
  assign net_40828 = seg_9_28_local_g1_2_40828;
  assign net_40831 = seg_9_28_local_g1_5_40831;
  assign net_40833 = seg_9_28_local_g1_7_40833;
  assign net_40836 = seg_9_28_local_g2_2_40836;
  assign net_40837 = seg_9_28_local_g2_3_40837;
  assign net_40839 = seg_9_28_local_g2_5_40839;
  assign net_40941 = seg_9_29_local_g0_0_40941;
  assign net_40950 = seg_9_29_local_g1_1_40950;
  assign net_40957 = seg_9_29_local_g2_0_40957;
  assign net_40960 = seg_9_29_local_g2_3_40960;
  assign net_40961 = seg_9_29_local_g2_4_40961;
  assign net_40962 = seg_9_29_local_g2_5_40962;
  assign net_40965 = seg_9_29_local_g3_0_40965;
  assign net_40970 = seg_9_29_local_g3_5_40970;
  assign net_41064 = seg_9_30_local_g0_0_41064;
  assign net_41068 = seg_9_30_local_g0_4_41068;
  assign net_41072 = seg_9_30_local_g1_0_41072;
  assign net_41077 = seg_9_30_local_g1_5_41077;
  assign net_41082 = seg_9_30_local_g2_2_41082;
  assign net_41083 = seg_9_30_local_g2_3_41083;
  assign net_41084 = seg_9_30_local_g2_4_41084;
  assign net_41094 = seg_9_30_local_g3_6_41094;
  assign net_41453 = seg_10_2_local_g0_2_41453;
  assign net_41454 = seg_10_2_local_g0_3_41454;
  assign net_41455 = seg_10_2_local_g0_4_41455;
  assign net_41457 = seg_10_2_local_g0_6_41457;
  assign net_41458 = seg_10_2_local_g0_7_41458;
  assign net_41462 = seg_10_2_local_g1_3_41462;
  assign net_41463 = seg_10_2_local_g1_4_41463;
  assign net_41465 = seg_10_2_local_g1_6_41465;
  assign net_41471 = seg_10_2_local_g2_4_41471;
  assign net_41477 = seg_10_2_local_g3_2_41477;
  assign net_41576 = seg_10_3_local_g0_2_41576;
  assign net_41585 = seg_10_3_local_g1_3_41585;
  assign net_41587 = seg_10_3_local_g1_5_41587;
  assign net_41588 = seg_10_3_local_g1_6_41588;
  assign net_41594 = seg_10_3_local_g2_4_41594;
  assign net_41600 = seg_10_3_local_g3_2_41600;
  assign net_41601 = seg_10_3_local_g3_3_41601;
  assign net_41605 = seg_10_3_local_g3_7_41605;
  assign net_42071 = seg_10_7_local_g0_5_42071;
  assign net_42082 = seg_10_7_local_g2_0_42082;
  assign net_42192 = seg_10_8_local_g0_3_42192;
  assign net_42194 = seg_10_8_local_g0_5_42194;
  assign net_42195 = seg_10_8_local_g0_6_42195;
  assign net_42196 = seg_10_8_local_g0_7_42196;
  assign net_42197 = seg_10_8_local_g1_0_42197;
  assign net_42200 = seg_10_8_local_g1_3_42200;
  assign net_42203 = seg_10_8_local_g1_6_42203;
  assign net_42205 = seg_10_8_local_g2_0_42205;
  assign net_42209 = seg_10_8_local_g2_4_42209;
  assign net_42210 = seg_10_8_local_g2_5_42210;
  assign net_42211 = seg_10_8_local_g2_6_42211;
  assign net_42212 = seg_10_8_local_g2_7_42212;
  assign net_42216 = seg_10_8_local_g3_3_42216;
  assign net_42220 = seg_10_8_local_g3_7_42220;
  assign net_42436 = seg_10_10_local_g0_1_42436;
  assign net_42441 = seg_10_10_local_g0_6_42441;
  assign net_42560 = seg_10_11_local_g0_2_42560;
  assign net_42563 = seg_10_11_local_g0_5_42563;
  assign net_42576 = seg_10_11_local_g2_2_42576;
  assign net_42578 = seg_10_11_local_g2_4_42578;
  assign net_42581 = seg_10_11_local_g2_7_42581;
  assign net_42586 = seg_10_11_local_g3_4_42586;
  assign net_42587 = seg_10_11_local_g3_5_42587;
  assign net_42681 = seg_10_12_local_g0_0_42681;
  assign net_42682 = seg_10_12_local_g0_1_42682;
  assign net_42684 = seg_10_12_local_g0_3_42684;
  assign net_42685 = seg_10_12_local_g0_4_42685;
  assign net_42686 = seg_10_12_local_g0_5_42686;
  assign net_42687 = seg_10_12_local_g0_6_42687;
  assign net_42689 = seg_10_12_local_g1_0_42689;
  assign net_42690 = seg_10_12_local_g1_1_42690;
  assign net_42692 = seg_10_12_local_g1_3_42692;
  assign net_42693 = seg_10_12_local_g1_4_42693;
  assign net_42696 = seg_10_12_local_g1_7_42696;
  assign net_42698 = seg_10_12_local_g2_1_42698;
  assign net_42699 = seg_10_12_local_g2_2_42699;
  assign net_42700 = seg_10_12_local_g2_3_42700;
  assign net_42702 = seg_10_12_local_g2_5_42702;
  assign net_42703 = seg_10_12_local_g2_6_42703;
  assign net_42708 = seg_10_12_local_g3_3_42708;
  assign net_42804 = seg_10_13_local_g0_0_42804;
  assign net_42805 = seg_10_13_local_g0_1_42805;
  assign net_42807 = seg_10_13_local_g0_3_42807;
  assign net_42808 = seg_10_13_local_g0_4_42808;
  assign net_42809 = seg_10_13_local_g0_5_42809;
  assign net_42810 = seg_10_13_local_g0_6_42810;
  assign net_42811 = seg_10_13_local_g0_7_42811;
  assign net_42812 = seg_10_13_local_g1_0_42812;
  assign net_42813 = seg_10_13_local_g1_1_42813;
  assign net_42815 = seg_10_13_local_g1_3_42815;
  assign net_42817 = seg_10_13_local_g1_5_42817;
  assign net_42822 = seg_10_13_local_g2_2_42822;
  assign net_42823 = seg_10_13_local_g2_3_42823;
  assign net_42828 = seg_10_13_local_g3_0_42828;
  assign net_42831 = seg_10_13_local_g3_3_42831;
  assign net_42832 = seg_10_13_local_g3_4_42832;
  assign net_42835 = seg_10_13_local_g3_7_42835;
  assign net_42927 = seg_10_14_local_g0_0_42927;
  assign net_42936 = seg_10_14_local_g1_1_42936;
  assign net_42938 = seg_10_14_local_g1_3_42938;
  assign net_42941 = seg_10_14_local_g1_6_42941;
  assign net_42942 = seg_10_14_local_g1_7_42942;
  assign net_42945 = seg_10_14_local_g2_2_42945;
  assign net_42947 = seg_10_14_local_g2_4_42947;
  assign net_42958 = seg_10_14_local_g3_7_42958;
  assign net_43052 = seg_10_15_local_g0_2_43052;
  assign net_43056 = seg_10_15_local_g0_6_43056;
  assign net_43074 = seg_10_15_local_g3_0_43074;
  assign net_43300 = seg_10_17_local_g0_4_43300;
  assign net_43302 = seg_10_17_local_g0_6_43302;
  assign net_43309 = seg_10_17_local_g1_5_43309;
  assign net_43311 = seg_10_17_local_g1_7_43311;
  assign net_43315 = seg_10_17_local_g2_3_43315;
  assign net_43321 = seg_10_17_local_g3_1_43321;
  assign net_43322 = seg_10_17_local_g3_2_43322;
  assign net_43325 = seg_10_17_local_g3_5_43325;
  assign net_43424 = seg_10_18_local_g0_5_43424;
  assign net_43430 = seg_10_18_local_g1_3_43430;
  assign net_43436 = seg_10_18_local_g2_1_43436;
  assign net_43437 = seg_10_18_local_g2_2_43437;
  assign net_43441 = seg_10_18_local_g2_6_43441;
  assign net_43443 = seg_10_18_local_g3_0_43443;
  assign net_43447 = seg_10_18_local_g3_4_43447;
  assign net_43450 = seg_10_18_local_g3_7_43450;
  assign net_43544 = seg_10_19_local_g0_2_43544;
  assign net_43548 = seg_10_19_local_g0_6_43548;
  assign net_43549 = seg_10_19_local_g0_7_43549;
  assign net_43550 = seg_10_19_local_g1_0_43550;
  assign net_43551 = seg_10_19_local_g1_1_43551;
  assign net_43554 = seg_10_19_local_g1_4_43554;
  assign net_43569 = seg_10_19_local_g3_3_43569;
  assign net_43571 = seg_10_19_local_g3_5_43571;
  assign net_43666 = seg_10_20_local_g0_1_43666;
  assign net_43668 = seg_10_20_local_g0_3_43668;
  assign net_43673 = seg_10_20_local_g1_0_43673;
  assign net_43691 = seg_10_20_local_g3_2_43691;
  assign net_44413 = seg_10_26_local_g1_2_44413;
  assign net_44430 = seg_10_26_local_g3_3_44430;
  assign net_44434 = seg_10_26_local_g3_7_44434;
  assign net_44529 = seg_10_27_local_g0_3_44529;
  assign net_44531 = seg_10_27_local_g0_5_44531;
  assign net_44532 = seg_10_27_local_g0_6_44532;
  assign net_44533 = seg_10_27_local_g0_7_44533;
  assign net_44537 = seg_10_27_local_g1_3_44537;
  assign net_44539 = seg_10_27_local_g1_5_44539;
  assign net_44541 = seg_10_27_local_g1_7_44541;
  assign net_44549 = seg_10_27_local_g2_7_44549;
  assign net_44553 = seg_10_27_local_g3_3_44553;
  assign net_44554 = seg_10_27_local_g3_4_44554;
  assign net_44653 = seg_10_28_local_g0_4_44653;
  assign net_44655 = seg_10_28_local_g0_6_44655;
  assign net_44656 = seg_10_28_local_g0_7_44656;
  assign net_44660 = seg_10_28_local_g1_3_44660;
  assign net_44663 = seg_10_28_local_g1_6_44663;
  assign net_44664 = seg_10_28_local_g1_7_44664;
  assign net_44670 = seg_10_28_local_g2_5_44670;
  assign net_44675 = seg_10_28_local_g3_2_44675;
  assign net_44676 = seg_10_28_local_g3_3_44676;
  assign net_44680 = seg_10_28_local_g3_7_44680;
  assign net_44773 = seg_10_29_local_g0_1_44773;
  assign net_44774 = seg_10_29_local_g0_2_44774;
  assign net_44783 = seg_10_29_local_g1_3_44783;
  assign net_44784 = seg_10_29_local_g1_4_44784;
  assign net_44788 = seg_10_29_local_g2_0_44788;
  assign net_44793 = seg_10_29_local_g2_5_44793;
  assign net_44803 = seg_10_29_local_g3_7_44803;
  assign net_44895 = seg_10_30_local_g0_0_44895;
  assign net_44897 = seg_10_30_local_g0_2_44897;
  assign net_44899 = seg_10_30_local_g0_4_44899;
  assign net_44900 = seg_10_30_local_g0_5_44900;
  assign net_44903 = seg_10_30_local_g1_0_44903;
  assign net_44905 = seg_10_30_local_g1_2_44905;
  assign net_44907 = seg_10_30_local_g1_4_44907;
  assign net_44908 = seg_10_30_local_g1_5_44908;
  assign net_44911 = seg_10_30_local_g2_0_44911;
  assign net_44913 = seg_10_30_local_g2_2_44913;
  assign net_44917 = seg_10_30_local_g2_6_44917;
  assign net_44922 = seg_10_30_local_g3_3_44922;
  assign net_44923 = seg_10_30_local_g3_4_44923;
  assign net_44925 = seg_10_30_local_g3_6_44925;
  assign net_44926 = seg_10_30_local_g3_7_44926;
  assign net_45907 = seg_11_7_local_g1_2_45907;
  assign net_45908 = seg_11_7_local_g1_3_45908;
  assign net_45911 = seg_11_7_local_g1_6_45911;
  assign net_45912 = seg_11_7_local_g1_7_45912;
  assign net_45921 = seg_11_7_local_g3_0_45921;
  assign net_45923 = seg_11_7_local_g3_2_45923;
  assign net_45924 = seg_11_7_local_g3_3_45924;
  assign net_46020 = seg_11_8_local_g0_0_46020;
  assign net_46021 = seg_11_8_local_g0_1_46021;
  assign net_46022 = seg_11_8_local_g0_2_46022;
  assign net_46023 = seg_11_8_local_g0_3_46023;
  assign net_46024 = seg_11_8_local_g0_4_46024;
  assign net_46028 = seg_11_8_local_g1_0_46028;
  assign net_46030 = seg_11_8_local_g1_2_46030;
  assign net_46034 = seg_11_8_local_g1_6_46034;
  assign net_46035 = seg_11_8_local_g1_7_46035;
  assign net_46037 = seg_11_8_local_g2_1_46037;
  assign net_46145 = seg_11_9_local_g0_2_46145;
  assign net_46146 = seg_11_9_local_g0_3_46146;
  assign net_46147 = seg_11_9_local_g0_4_46147;
  assign net_46148 = seg_11_9_local_g0_5_46148;
  assign net_46149 = seg_11_9_local_g0_6_46149;
  assign net_46150 = seg_11_9_local_g0_7_46150;
  assign net_46154 = seg_11_9_local_g1_3_46154;
  assign net_46155 = seg_11_9_local_g1_4_46155;
  assign net_46156 = seg_11_9_local_g1_5_46156;
  assign net_46157 = seg_11_9_local_g1_6_46157;
  assign net_46158 = seg_11_9_local_g1_7_46158;
  assign net_46165 = seg_11_9_local_g2_6_46165;
  assign net_46167 = seg_11_9_local_g3_0_46167;
  assign net_46268 = seg_11_10_local_g0_2_46268;
  assign net_46269 = seg_11_10_local_g0_3_46269;
  assign net_46271 = seg_11_10_local_g0_5_46271;
  assign net_46273 = seg_11_10_local_g0_7_46273;
  assign net_46276 = seg_11_10_local_g1_2_46276;
  assign net_46277 = seg_11_10_local_g1_3_46277;
  assign net_46279 = seg_11_10_local_g1_5_46279;
  assign net_46286 = seg_11_10_local_g2_4_46286;
  assign net_46292 = seg_11_10_local_g3_2_46292;
  assign net_46294 = seg_11_10_local_g3_4_46294;
  assign net_46297 = seg_11_10_local_g3_7_46297;
  assign net_46407 = seg_11_11_local_g2_2_46407;
  assign net_46419 = seg_11_11_local_g3_6_46419;
  assign net_46513 = seg_11_12_local_g0_1_46513;
  assign net_46514 = seg_11_12_local_g0_2_46514;
  assign net_46517 = seg_11_12_local_g0_5_46517;
  assign net_46519 = seg_11_12_local_g0_7_46519;
  assign net_46525 = seg_11_12_local_g1_5_46525;
  assign net_46529 = seg_11_12_local_g2_1_46529;
  assign net_46532 = seg_11_12_local_g2_4_46532;
  assign net_46533 = seg_11_12_local_g2_5_46533;
  assign net_46534 = seg_11_12_local_g2_6_46534;
  assign net_46535 = seg_11_12_local_g2_7_46535;
  assign net_46537 = seg_11_12_local_g3_1_46537;
  assign net_46639 = seg_11_13_local_g0_4_46639;
  assign net_46640 = seg_11_13_local_g0_5_46640;
  assign net_46641 = seg_11_13_local_g0_6_46641;
  assign net_46642 = seg_11_13_local_g0_7_46642;
  assign net_46644 = seg_11_13_local_g1_1_46644;
  assign net_46645 = seg_11_13_local_g1_2_46645;
  assign net_46646 = seg_11_13_local_g1_3_46646;
  assign net_46647 = seg_11_13_local_g1_4_46647;
  assign net_46648 = seg_11_13_local_g1_5_46648;
  assign net_46650 = seg_11_13_local_g1_7_46650;
  assign net_46652 = seg_11_13_local_g2_1_46652;
  assign net_46653 = seg_11_13_local_g2_2_46653;
  assign net_46656 = seg_11_13_local_g2_5_46656;
  assign net_46658 = seg_11_13_local_g2_7_46658;
  assign net_46663 = seg_11_13_local_g3_4_46663;
  assign net_46665 = seg_11_13_local_g3_6_46665;
  assign net_46758 = seg_11_14_local_g0_0_46758;
  assign net_46760 = seg_11_14_local_g0_2_46760;
  assign net_46762 = seg_11_14_local_g0_4_46762;
  assign net_46764 = seg_11_14_local_g0_6_46764;
  assign net_46765 = seg_11_14_local_g0_7_46765;
  assign net_46768 = seg_11_14_local_g1_2_46768;
  assign net_46769 = seg_11_14_local_g1_3_46769;
  assign net_46773 = seg_11_14_local_g1_7_46773;
  assign net_46774 = seg_11_14_local_g2_0_46774;
  assign net_46776 = seg_11_14_local_g2_2_46776;
  assign net_46780 = seg_11_14_local_g2_6_46780;
  assign net_46784 = seg_11_14_local_g3_2_46784;
  assign net_46884 = seg_11_15_local_g0_3_46884;
  assign net_46892 = seg_11_15_local_g1_3_46892;
  assign net_46894 = seg_11_15_local_g1_5_46894;
  assign net_46898 = seg_11_15_local_g2_1_46898;
  assign net_46905 = seg_11_15_local_g3_0_46905;
  assign net_47006 = seg_11_16_local_g0_2_47006;
  assign net_47009 = seg_11_16_local_g0_5_47009;
  assign net_47128 = seg_11_17_local_g0_1_47128;
  assign net_47148 = seg_11_17_local_g2_5_47148;
  assign net_47252 = seg_11_18_local_g0_2_47252;
  assign net_47258 = seg_11_18_local_g1_0_47258;
  assign net_47268 = seg_11_18_local_g2_2_47268;
  assign net_47269 = seg_11_18_local_g2_3_47269;
  assign net_47271 = seg_11_18_local_g2_5_47271;
  assign net_47272 = seg_11_18_local_g2_6_47272;
  assign net_47274 = seg_11_18_local_g3_0_47274;
  assign net_47275 = seg_11_18_local_g3_1_47275;
  assign net_47276 = seg_11_18_local_g3_2_47276;
  assign net_47279 = seg_11_18_local_g3_5_47279;
  assign net_47374 = seg_11_19_local_g0_1_47374;
  assign net_47377 = seg_11_19_local_g0_4_47377;
  assign net_47382 = seg_11_19_local_g1_1_47382;
  assign net_47385 = seg_11_19_local_g1_4_47385;
  assign net_47391 = seg_11_19_local_g2_2_47391;
  assign net_47397 = seg_11_19_local_g3_0_47397;
  assign net_47403 = seg_11_19_local_g3_6_47403;
  assign net_47498 = seg_11_20_local_g0_2_47498;
  assign net_47505 = seg_11_20_local_g1_1_47505;
  assign net_47516 = seg_11_20_local_g2_4_47516;
  assign net_47883 = seg_11_23_local_g2_2_47883;
  assign net_47892 = seg_11_23_local_g3_3_47892;
  assign net_48606 = seg_11_29_local_g0_3_48606;
  assign net_48616 = seg_11_29_local_g1_5_48616;
  assign net_48737 = seg_11_30_local_g1_3_48737;
  assign net_48738 = seg_11_30_local_g1_4_48738;
  assign net_48742 = seg_11_30_local_g2_0_48742;
  assign net_48747 = seg_11_30_local_g2_5_48747;
  assign net_49862 = seg_12_8_local_g1_3_49862;
  assign net_49866 = seg_12_8_local_g1_7_49866;
  assign net_49872 = seg_12_8_local_g2_5_49872;
  assign net_49875 = seg_12_8_local_g3_0_49875;
  assign net_49876 = seg_12_8_local_g3_1_49876;
  assign net_49880 = seg_12_8_local_g3_5_49880;
  assign net_5 = seg_23_9_glb_netwk_0_5;
  assign net_50220 = seg_12_11_local_g0_0_50220;
  assign net_50223 = seg_12_11_local_g0_3_50223;
  assign net_50226 = seg_12_11_local_g0_6_50226;
  assign net_50227 = seg_12_11_local_g0_7_50227;
  assign net_50229 = seg_12_11_local_g1_1_50229;
  assign net_50230 = seg_12_11_local_g1_2_50230;
  assign net_50234 = seg_12_11_local_g1_6_50234;
  assign net_50239 = seg_12_11_local_g2_3_50239;
  assign net_50240 = seg_12_11_local_g2_4_50240;
  assign net_50247 = seg_12_11_local_g3_3_50247;
  assign net_50343 = seg_12_12_local_g0_0_50343;
  assign net_50344 = seg_12_12_local_g0_1_50344;
  assign net_50345 = seg_12_12_local_g0_2_50345;
  assign net_50346 = seg_12_12_local_g0_3_50346;
  assign net_50347 = seg_12_12_local_g0_4_50347;
  assign net_50348 = seg_12_12_local_g0_5_50348;
  assign net_50349 = seg_12_12_local_g0_6_50349;
  assign net_50351 = seg_12_12_local_g1_0_50351;
  assign net_50353 = seg_12_12_local_g1_2_50353;
  assign net_50354 = seg_12_12_local_g1_3_50354;
  assign net_50355 = seg_12_12_local_g1_4_50355;
  assign net_50356 = seg_12_12_local_g1_5_50356;
  assign net_50359 = seg_12_12_local_g2_0_50359;
  assign net_50360 = seg_12_12_local_g2_1_50360;
  assign net_50361 = seg_12_12_local_g2_2_50361;
  assign net_50370 = seg_12_12_local_g3_3_50370;
  assign net_50371 = seg_12_12_local_g3_4_50371;
  assign net_50466 = seg_12_13_local_g0_0_50466;
  assign net_50467 = seg_12_13_local_g0_1_50467;
  assign net_50468 = seg_12_13_local_g0_2_50468;
  assign net_50469 = seg_12_13_local_g0_3_50469;
  assign net_50471 = seg_12_13_local_g0_5_50471;
  assign net_50474 = seg_12_13_local_g1_0_50474;
  assign net_50475 = seg_12_13_local_g1_1_50475;
  assign net_50477 = seg_12_13_local_g1_3_50477;
  assign net_50478 = seg_12_13_local_g1_4_50478;
  assign net_50479 = seg_12_13_local_g1_5_50479;
  assign net_50481 = seg_12_13_local_g1_7_50481;
  assign net_50483 = seg_12_13_local_g2_1_50483;
  assign net_50484 = seg_12_13_local_g2_2_50484;
  assign net_50485 = seg_12_13_local_g2_3_50485;
  assign net_50492 = seg_12_13_local_g3_2_50492;
  assign net_50493 = seg_12_13_local_g3_3_50493;
  assign net_50495 = seg_12_13_local_g3_5_50495;
  assign net_50593 = seg_12_14_local_g0_4_50593;
  assign net_50597 = seg_12_14_local_g1_0_50597;
  assign net_50598 = seg_12_14_local_g1_1_50598;
  assign net_50599 = seg_12_14_local_g1_2_50599;
  assign net_50600 = seg_12_14_local_g1_3_50600;
  assign net_50601 = seg_12_14_local_g1_4_50601;
  assign net_50602 = seg_12_14_local_g1_5_50602;
  assign net_50603 = seg_12_14_local_g1_6_50603;
  assign net_50609 = seg_12_14_local_g2_4_50609;
  assign net_50613 = seg_12_14_local_g3_0_50613;
  assign net_50615 = seg_12_14_local_g3_2_50615;
  assign net_50616 = seg_12_14_local_g3_3_50616;
  assign net_50617 = seg_12_14_local_g3_4_50617;
  assign net_50620 = seg_12_14_local_g3_7_50620;
  assign net_50712 = seg_12_15_local_g0_0_50712;
  assign net_50713 = seg_12_15_local_g0_1_50713;
  assign net_50716 = seg_12_15_local_g0_4_50716;
  assign net_50718 = seg_12_15_local_g0_6_50718;
  assign net_50722 = seg_12_15_local_g1_2_50722;
  assign net_50724 = seg_12_15_local_g1_4_50724;
  assign net_50726 = seg_12_15_local_g1_6_50726;
  assign net_50728 = seg_12_15_local_g2_0_50728;
  assign net_50735 = seg_12_15_local_g2_7_50735;
  assign net_50740 = seg_12_15_local_g3_4_50740;
  assign net_50743 = seg_12_15_local_g3_7_50743;
  assign net_50835 = seg_12_16_local_g0_0_50835;
  assign net_50836 = seg_12_16_local_g0_1_50836;
  assign net_50854 = seg_12_16_local_g2_3_50854;
  assign net_50861 = seg_12_16_local_g3_2_50861;
  assign net_50862 = seg_12_16_local_g3_3_50862;
  assign net_50865 = seg_12_16_local_g3_6_50865;
  assign net_50960 = seg_12_17_local_g0_2_50960;
  assign net_50962 = seg_12_17_local_g0_4_50962;
  assign net_50963 = seg_12_17_local_g0_5_50963;
  assign net_50967 = seg_12_17_local_g1_1_50967;
  assign net_50971 = seg_12_17_local_g1_5_50971;
  assign net_50980 = seg_12_17_local_g2_6_50980;
  assign net_51082 = seg_12_18_local_g0_1_51082;
  assign net_51085 = seg_12_18_local_g0_4_51085;
  assign net_51086 = seg_12_18_local_g0_5_51086;
  assign net_51088 = seg_12_18_local_g0_7_51088;
  assign net_51095 = seg_12_18_local_g1_6_51095;
  assign net_51099 = seg_12_18_local_g2_2_51099;
  assign net_51101 = seg_12_18_local_g2_4_51101;
  assign net_51103 = seg_12_18_local_g2_6_51103;
  assign net_51105 = seg_12_18_local_g3_0_51105;
  assign net_51106 = seg_12_18_local_g3_1_51106;
  assign net_51210 = seg_12_19_local_g0_6_51210;
  assign net_51213 = seg_12_19_local_g1_1_51213;
  assign net_51214 = seg_12_19_local_g1_2_51214;
  assign net_51215 = seg_12_19_local_g1_3_51215;
  assign net_51216 = seg_12_19_local_g1_4_51216;
  assign net_51220 = seg_12_19_local_g2_0_51220;
  assign net_51222 = seg_12_19_local_g2_2_51222;
  assign net_51228 = seg_12_19_local_g3_0_51228;
  assign net_51231 = seg_12_19_local_g3_3_51231;
  assign net_51235 = seg_12_19_local_g3_7_51235;
  assign net_51343 = seg_12_20_local_g2_0_51343;
  assign net_51452 = seg_12_21_local_g0_2_51452;
  assign net_51456 = seg_12_21_local_g0_6_51456;
  assign net_51460 = seg_12_21_local_g1_2_51460;
  assign net_51461 = seg_12_21_local_g1_3_51461;
  assign net_51470 = seg_12_21_local_g2_4_51470;
  assign net_51471 = seg_12_21_local_g2_5_51471;
  assign net_51473 = seg_12_21_local_g2_7_51473;
  assign net_51477 = seg_12_21_local_g3_3_51477;
  assign net_51719 = seg_12_23_local_g2_7_51719;
  assign net_52195 = seg_12_27_local_g0_7_52195;
  assign net_52197 = seg_12_27_local_g1_1_52197;
  assign net_52199 = seg_12_27_local_g1_3_52199;
  assign net_52206 = seg_12_27_local_g2_2_52206;
  assign net_52207 = seg_12_27_local_g2_3_52207;
  assign net_52208 = seg_12_27_local_g2_4_52208;
  assign net_52209 = seg_12_27_local_g2_5_52209;
  assign net_52211 = seg_12_27_local_g2_7_52211;
  assign net_52215 = seg_12_27_local_g3_3_52215;
  assign net_52218 = seg_12_27_local_g3_6_52218;
  assign net_52313 = seg_12_28_local_g0_2_52313;
  assign net_52320 = seg_12_28_local_g1_1_52320;
  assign net_52321 = seg_12_28_local_g1_2_52321;
  assign net_52322 = seg_12_28_local_g1_3_52322;
  assign net_52336 = seg_12_28_local_g3_1_52336;
  assign net_53073 = seg_13_3_local_g0_6_53073;
  assign net_53074 = seg_13_3_local_g0_7_53074;
  assign net_53078 = seg_13_3_local_g1_3_53078;
  assign net_53092 = seg_13_3_local_g3_1_53092;
  assign net_53095 = seg_13_3_local_g3_4_53095;
  assign net_53098 = seg_13_3_local_g3_7_53098;
  assign net_53194 = seg_13_4_local_g0_4_53194;
  assign net_53198 = seg_13_4_local_g1_0_53198;
  assign net_53204 = seg_13_4_local_g1_6_53204;
  assign net_53208 = seg_13_4_local_g2_2_53208;
  assign net_53210 = seg_13_4_local_g2_4_53210;
  assign net_53211 = seg_13_4_local_g2_5_53211;
  assign net_53213 = seg_13_4_local_g2_7_53213;
  assign net_53214 = seg_13_4_local_g3_0_53214;
  assign net_53215 = seg_13_4_local_g3_1_53215;
  assign net_53221 = seg_13_4_local_g3_7_53221;
  assign net_53682 = seg_13_8_local_g0_0_53682;
  assign net_53683 = seg_13_8_local_g0_1_53683;
  assign net_53687 = seg_13_8_local_g0_5_53687;
  assign net_53688 = seg_13_8_local_g0_6_53688;
  assign net_53690 = seg_13_8_local_g1_0_53690;
  assign net_53696 = seg_13_8_local_g1_6_53696;
  assign net_53712 = seg_13_8_local_g3_6_53712;
  assign net_53713 = seg_13_8_local_g3_7_53713;
  assign net_53807 = seg_13_9_local_g0_2_53807;
  assign net_53809 = seg_13_9_local_g0_4_53809;
  assign net_53814 = seg_13_9_local_g1_1_53814;
  assign net_53815 = seg_13_9_local_g1_2_53815;
  assign net_53817 = seg_13_9_local_g1_4_53817;
  assign net_53818 = seg_13_9_local_g1_5_53818;
  assign net_53819 = seg_13_9_local_g1_6_53819;
  assign net_53820 = seg_13_9_local_g1_7_53820;
  assign net_53823 = seg_13_9_local_g2_2_53823;
  assign net_53825 = seg_13_9_local_g2_4_53825;
  assign net_53827 = seg_13_9_local_g2_6_53827;
  assign net_53831 = seg_13_9_local_g3_2_53831;
  assign net_53832 = seg_13_9_local_g3_3_53832;
  assign net_53834 = seg_13_9_local_g3_5_53834;
  assign net_53836 = seg_13_9_local_g3_7_53836;
  assign net_54064 = seg_13_11_local_g1_5_54064;
  assign net_54069 = seg_13_11_local_g2_2_54069;
  assign net_54081 = seg_13_11_local_g3_6_54081;
  assign net_54175 = seg_13_12_local_g0_1_54175;
  assign net_54176 = seg_13_12_local_g0_2_54176;
  assign net_54177 = seg_13_12_local_g0_3_54177;
  assign net_54178 = seg_13_12_local_g0_4_54178;
  assign net_54179 = seg_13_12_local_g0_5_54179;
  assign net_54186 = seg_13_12_local_g1_4_54186;
  assign net_54187 = seg_13_12_local_g1_5_54187;
  assign net_54188 = seg_13_12_local_g1_6_54188;
  assign net_54189 = seg_13_12_local_g1_7_54189;
  assign net_54190 = seg_13_12_local_g2_0_54190;
  assign net_54191 = seg_13_12_local_g2_1_54191;
  assign net_54193 = seg_13_12_local_g2_3_54193;
  assign net_54195 = seg_13_12_local_g2_5_54195;
  assign net_54202 = seg_13_12_local_g3_4_54202;
  assign net_54205 = seg_13_12_local_g3_7_54205;
  assign net_54297 = seg_13_13_local_g0_0_54297;
  assign net_54299 = seg_13_13_local_g0_2_54299;
  assign net_54300 = seg_13_13_local_g0_3_54300;
  assign net_54302 = seg_13_13_local_g0_5_54302;
  assign net_54305 = seg_13_13_local_g1_0_54305;
  assign net_54308 = seg_13_13_local_g1_3_54308;
  assign net_54309 = seg_13_13_local_g1_4_54309;
  assign net_54310 = seg_13_13_local_g1_5_54310;
  assign net_54312 = seg_13_13_local_g1_7_54312;
  assign net_54316 = seg_13_13_local_g2_3_54316;
  assign net_54318 = seg_13_13_local_g2_5_54318;
  assign net_54319 = seg_13_13_local_g2_6_54319;
  assign net_54323 = seg_13_13_local_g3_2_54323;
  assign net_54325 = seg_13_13_local_g3_4_54325;
  assign net_54326 = seg_13_13_local_g3_5_54326;
  assign net_54328 = seg_13_13_local_g3_7_54328;
  assign net_54426 = seg_13_14_local_g0_6_54426;
  assign net_54427 = seg_13_14_local_g0_7_54427;
  assign net_54428 = seg_13_14_local_g1_0_54428;
  assign net_54431 = seg_13_14_local_g1_3_54431;
  assign net_54433 = seg_13_14_local_g1_5_54433;
  assign net_54434 = seg_13_14_local_g1_6_54434;
  assign net_54435 = seg_13_14_local_g1_7_54435;
  assign net_54437 = seg_13_14_local_g2_1_54437;
  assign net_54442 = seg_13_14_local_g2_6_54442;
  assign net_54444 = seg_13_14_local_g3_0_54444;
  assign net_54446 = seg_13_14_local_g3_2_54446;
  assign net_54447 = seg_13_14_local_g3_3_54447;
  assign net_54449 = seg_13_14_local_g3_5_54449;
  assign net_54450 = seg_13_14_local_g3_6_54450;
  assign net_54451 = seg_13_14_local_g3_7_54451;
  assign net_54545 = seg_13_15_local_g0_2_54545;
  assign net_54548 = seg_13_15_local_g0_5_54548;
  assign net_54553 = seg_13_15_local_g1_2_54553;
  assign net_54555 = seg_13_15_local_g1_4_54555;
  assign net_54559 = seg_13_15_local_g2_0_54559;
  assign net_54560 = seg_13_15_local_g2_1_54560;
  assign net_54561 = seg_13_15_local_g2_2_54561;
  assign net_54562 = seg_13_15_local_g2_3_54562;
  assign net_54564 = seg_13_15_local_g2_5_54564;
  assign net_54565 = seg_13_15_local_g2_6_54565;
  assign net_54569 = seg_13_15_local_g3_2_54569;
  assign net_54570 = seg_13_15_local_g3_3_54570;
  assign net_54572 = seg_13_15_local_g3_5_54572;
  assign net_54573 = seg_13_15_local_g3_6_54573;
  assign net_54668 = seg_13_16_local_g0_2_54668;
  assign net_54670 = seg_13_16_local_g0_4_54670;
  assign net_54672 = seg_13_16_local_g0_6_54672;
  assign net_54677 = seg_13_16_local_g1_3_54677;
  assign net_54680 = seg_13_16_local_g1_6_54680;
  assign net_54682 = seg_13_16_local_g2_0_54682;
  assign net_54685 = seg_13_16_local_g2_3_54685;
  assign net_54686 = seg_13_16_local_g2_4_54686;
  assign net_54687 = seg_13_16_local_g2_5_54687;
  assign net_54689 = seg_13_16_local_g2_7_54689;
  assign net_54690 = seg_13_16_local_g3_0_54690;
  assign net_54692 = seg_13_16_local_g3_2_54692;
  assign net_54693 = seg_13_16_local_g3_3_54693;
  assign net_54694 = seg_13_16_local_g3_4_54694;
  assign net_54695 = seg_13_16_local_g3_5_54695;
  assign net_54696 = seg_13_16_local_g3_6_54696;
  assign net_54697 = seg_13_16_local_g3_7_54697;
  assign net_54789 = seg_13_17_local_g0_0_54789;
  assign net_54792 = seg_13_17_local_g0_3_54792;
  assign net_54793 = seg_13_17_local_g0_4_54793;
  assign net_54795 = seg_13_17_local_g0_6_54795;
  assign net_54797 = seg_13_17_local_g1_0_54797;
  assign net_54801 = seg_13_17_local_g1_4_54801;
  assign net_54803 = seg_13_17_local_g1_6_54803;
  assign net_54805 = seg_13_17_local_g2_0_54805;
  assign net_54806 = seg_13_17_local_g2_1_54806;
  assign net_54808 = seg_13_17_local_g2_3_54808;
  assign net_54811 = seg_13_17_local_g2_6_54811;
  assign net_54812 = seg_13_17_local_g2_7_54812;
  assign net_54814 = seg_13_17_local_g3_1_54814;
  assign net_54815 = seg_13_17_local_g3_2_54815;
  assign net_54816 = seg_13_17_local_g3_3_54816;
  assign net_54818 = seg_13_17_local_g3_5_54818;
  assign net_54820 = seg_13_17_local_g3_7_54820;
  assign net_54912 = seg_13_18_local_g0_0_54912;
  assign net_54933 = seg_13_18_local_g2_5_54933;
  assign net_54943 = seg_13_18_local_g3_7_54943;
  assign net_55042 = seg_13_19_local_g0_7_55042;
  assign net_55043 = seg_13_19_local_g1_0_55043;
  assign net_55049 = seg_13_19_local_g1_6_55049;
  assign net_55050 = seg_13_19_local_g1_7_55050;
  assign net_55052 = seg_13_19_local_g2_1_55052;
  assign net_55053 = seg_13_19_local_g2_2_55053;
  assign net_55055 = seg_13_19_local_g2_4_55055;
  assign net_55056 = seg_13_19_local_g2_5_55056;
  assign net_55057 = seg_13_19_local_g2_6_55057;
  assign net_55058 = seg_13_19_local_g2_7_55058;
  assign net_55062 = seg_13_19_local_g3_3_55062;
  assign net_55063 = seg_13_19_local_g3_4_55063;
  assign net_55064 = seg_13_19_local_g3_5_55064;
  assign net_55066 = seg_13_19_local_g3_7_55066;
  assign net_55169 = seg_13_20_local_g1_3_55169;
  assign net_55171 = seg_13_20_local_g1_5_55171;
  assign net_55172 = seg_13_20_local_g1_6_55172;
  assign net_55175 = seg_13_20_local_g2_1_55175;
  assign net_55176 = seg_13_20_local_g2_2_55176;
  assign net_55178 = seg_13_20_local_g2_4_55178;
  assign net_55181 = seg_13_20_local_g2_7_55181;
  assign net_55182 = seg_13_20_local_g3_0_55182;
  assign net_55183 = seg_13_20_local_g3_1_55183;
  assign net_55186 = seg_13_20_local_g3_4_55186;
  assign net_55187 = seg_13_20_local_g3_5_55187;
  assign net_55189 = seg_13_20_local_g3_7_55189;
  assign net_55309 = seg_13_21_local_g3_4_55309;
  assign net_55405 = seg_13_22_local_g0_1_55405;
  assign net_55417 = seg_13_22_local_g1_5_55417;
  assign net_55418 = seg_13_22_local_g1_6_55418;
  assign net_55422 = seg_13_22_local_g2_2_55422;
  assign net_55423 = seg_13_22_local_g2_3_55423;
  assign net_55433 = seg_13_22_local_g3_5_55433;
  assign net_56021 = seg_13_27_local_g0_2_56021;
  assign net_56024 = seg_13_27_local_g0_5_56024;
  assign net_56025 = seg_13_27_local_g0_6_56025;
  assign net_56026 = seg_13_27_local_g0_7_56026;
  assign net_56030 = seg_13_27_local_g1_3_56030;
  assign net_56031 = seg_13_27_local_g1_4_56031;
  assign net_56034 = seg_13_27_local_g1_7_56034;
  assign net_56036 = seg_13_27_local_g2_1_56036;
  assign net_56037 = seg_13_27_local_g2_2_56037;
  assign net_56040 = seg_13_27_local_g2_5_56040;
  assign net_56047 = seg_13_27_local_g3_4_56047;
  assign net_56534 = seg_13_31_local_g1_2_56534;
  assign net_56535 = seg_13_31_local_g1_3_56535;
  assign net_56776 = seg_14_2_local_g0_2_56776;
  assign net_56777 = seg_14_2_local_g0_3_56777;
  assign net_56780 = seg_14_2_local_g0_6_56780;
  assign net_56785 = seg_14_2_local_g1_3_56785;
  assign net_56790 = seg_14_2_local_g2_0_56790;
  assign net_56793 = seg_14_2_local_g2_3_56793;
  assign net_56800 = seg_14_2_local_g3_2_56800;
  assign net_56805 = seg_14_2_local_g3_7_56805;
  assign net_56897 = seg_14_3_local_g0_0_56897;
  assign net_56898 = seg_14_3_local_g0_1_56898;
  assign net_56899 = seg_14_3_local_g0_2_56899;
  assign net_56904 = seg_14_3_local_g0_7_56904;
  assign net_56905 = seg_14_3_local_g1_0_56905;
  assign net_56906 = seg_14_3_local_g1_1_56906;
  assign net_56908 = seg_14_3_local_g1_3_56908;
  assign net_56909 = seg_14_3_local_g1_4_56909;
  assign net_56911 = seg_14_3_local_g1_6_56911;
  assign net_56912 = seg_14_3_local_g1_7_56912;
  assign net_56914 = seg_14_3_local_g2_1_56914;
  assign net_56915 = seg_14_3_local_g2_2_56915;
  assign net_56916 = seg_14_3_local_g2_3_56916;
  assign net_56917 = seg_14_3_local_g2_4_56917;
  assign net_56920 = seg_14_3_local_g2_7_56920;
  assign net_56921 = seg_14_3_local_g3_0_56921;
  assign net_56924 = seg_14_3_local_g3_3_56924;
  assign net_56928 = seg_14_3_local_g3_7_56928;
  assign net_57023 = seg_14_4_local_g0_3_57023;
  assign net_57027 = seg_14_4_local_g0_7_57027;
  assign net_57028 = seg_14_4_local_g1_0_57028;
  assign net_57030 = seg_14_4_local_g1_2_57030;
  assign net_57034 = seg_14_4_local_g1_6_57034;
  assign net_57038 = seg_14_4_local_g2_2_57038;
  assign net_57041 = seg_14_4_local_g2_5_57041;
  assign net_57044 = seg_14_4_local_g3_0_57044;
  assign net_57046 = seg_14_4_local_g3_2_57046;
  assign net_57049 = seg_14_4_local_g3_5_57049;
  assign net_57051 = seg_14_4_local_g3_7_57051;
  assign net_57391 = seg_14_7_local_g0_2_57391;
  assign net_57403 = seg_14_7_local_g1_6_57403;
  assign net_57410 = seg_14_7_local_g2_5_57410;
  assign net_57412 = seg_14_7_local_g2_7_57412;
  assign net_57414 = seg_14_7_local_g3_1_57414;
  assign net_57415 = seg_14_7_local_g3_2_57415;
  assign net_57418 = seg_14_7_local_g3_5_57418;
  assign net_57515 = seg_14_8_local_g0_3_57515;
  assign net_57518 = seg_14_8_local_g0_6_57518;
  assign net_57523 = seg_14_8_local_g1_3_57523;
  assign net_57526 = seg_14_8_local_g1_6_57526;
  assign net_57527 = seg_14_8_local_g1_7_57527;
  assign net_57528 = seg_14_8_local_g2_0_57528;
  assign net_57529 = seg_14_8_local_g2_1_57529;
  assign net_57535 = seg_14_8_local_g2_7_57535;
  assign net_57536 = seg_14_8_local_g3_0_57536;
  assign net_57539 = seg_14_8_local_g3_3_57539;
  assign net_57541 = seg_14_8_local_g3_5_57541;
  assign net_57543 = seg_14_8_local_g3_7_57543;
  assign net_57635 = seg_14_9_local_g0_0_57635;
  assign net_57636 = seg_14_9_local_g0_1_57636;
  assign net_57640 = seg_14_9_local_g0_5_57640;
  assign net_57641 = seg_14_9_local_g0_6_57641;
  assign net_57642 = seg_14_9_local_g0_7_57642;
  assign net_57643 = seg_14_9_local_g1_0_57643;
  assign net_57647 = seg_14_9_local_g1_4_57647;
  assign net_57649 = seg_14_9_local_g1_6_57649;
  assign net_57652 = seg_14_9_local_g2_1_57652;
  assign net_57660 = seg_14_9_local_g3_1_57660;
  assign net_57763 = seg_14_10_local_g0_5_57763;
  assign net_57764 = seg_14_10_local_g0_6_57764;
  assign net_57776 = seg_14_10_local_g2_2_57776;
  assign net_57779 = seg_14_10_local_g2_5_57779;
  assign net_57884 = seg_14_11_local_g0_3_57884;
  assign net_57885 = seg_14_11_local_g0_4_57885;
  assign net_57887 = seg_14_11_local_g0_6_57887;
  assign net_57888 = seg_14_11_local_g0_7_57888;
  assign net_57890 = seg_14_11_local_g1_1_57890;
  assign net_57893 = seg_14_11_local_g1_4_57893;
  assign net_57897 = seg_14_11_local_g2_0_57897;
  assign net_57899 = seg_14_11_local_g2_2_57899;
  assign net_57900 = seg_14_11_local_g2_3_57900;
  assign net_57902 = seg_14_11_local_g2_5_57902;
  assign net_57903 = seg_14_11_local_g2_6_57903;
  assign net_58006 = seg_14_12_local_g0_2_58006;
  assign net_58007 = seg_14_12_local_g0_3_58007;
  assign net_58012 = seg_14_12_local_g1_0_58012;
  assign net_58013 = seg_14_12_local_g1_1_58013;
  assign net_58014 = seg_14_12_local_g1_2_58014;
  assign net_58015 = seg_14_12_local_g1_3_58015;
  assign net_58018 = seg_14_12_local_g1_6_58018;
  assign net_58019 = seg_14_12_local_g1_7_58019;
  assign net_58021 = seg_14_12_local_g2_1_58021;
  assign net_58023 = seg_14_12_local_g2_3_58023;
  assign net_58024 = seg_14_12_local_g2_4_58024;
  assign net_58026 = seg_14_12_local_g2_6_58026;
  assign net_58027 = seg_14_12_local_g2_7_58027;
  assign net_58031 = seg_14_12_local_g3_3_58031;
  assign net_58034 = seg_14_12_local_g3_6_58034;
  assign net_58035 = seg_14_12_local_g3_7_58035;
  assign net_58128 = seg_14_13_local_g0_1_58128;
  assign net_58129 = seg_14_13_local_g0_2_58129;
  assign net_58130 = seg_14_13_local_g0_3_58130;
  assign net_58133 = seg_14_13_local_g0_6_58133;
  assign net_58134 = seg_14_13_local_g0_7_58134;
  assign net_58135 = seg_14_13_local_g1_0_58135;
  assign net_58136 = seg_14_13_local_g1_1_58136;
  assign net_58137 = seg_14_13_local_g1_2_58137;
  assign net_58138 = seg_14_13_local_g1_3_58138;
  assign net_58140 = seg_14_13_local_g1_5_58140;
  assign net_58141 = seg_14_13_local_g1_6_58141;
  assign net_58142 = seg_14_13_local_g1_7_58142;
  assign net_58144 = seg_14_13_local_g2_1_58144;
  assign net_58145 = seg_14_13_local_g2_2_58145;
  assign net_58147 = seg_14_13_local_g2_4_58147;
  assign net_58148 = seg_14_13_local_g2_5_58148;
  assign net_58149 = seg_14_13_local_g2_6_58149;
  assign net_58150 = seg_14_13_local_g2_7_58150;
  assign net_58151 = seg_14_13_local_g3_0_58151;
  assign net_58152 = seg_14_13_local_g3_1_58152;
  assign net_58154 = seg_14_13_local_g3_3_58154;
  assign net_58155 = seg_14_13_local_g3_4_58155;
  assign net_58156 = seg_14_13_local_g3_5_58156;
  assign net_58157 = seg_14_13_local_g3_6_58157;
  assign net_58158 = seg_14_13_local_g3_7_58158;
  assign net_58258 = seg_14_14_local_g1_0_58258;
  assign net_58260 = seg_14_14_local_g1_2_58260;
  assign net_58261 = seg_14_14_local_g1_3_58261;
  assign net_58262 = seg_14_14_local_g1_4_58262;
  assign net_58263 = seg_14_14_local_g1_5_58263;
  assign net_58264 = seg_14_14_local_g1_6_58264;
  assign net_58270 = seg_14_14_local_g2_4_58270;
  assign net_58272 = seg_14_14_local_g2_6_58272;
  assign net_58273 = seg_14_14_local_g2_7_58273;
  assign net_58274 = seg_14_14_local_g3_0_58274;
  assign net_58276 = seg_14_14_local_g3_2_58276;
  assign net_58277 = seg_14_14_local_g3_3_58277;
  assign net_58279 = seg_14_14_local_g3_5_58279;
  assign net_58280 = seg_14_14_local_g3_6_58280;
  assign net_58281 = seg_14_14_local_g3_7_58281;
  assign net_58382 = seg_14_15_local_g1_1_58382;
  assign net_58383 = seg_14_15_local_g1_2_58383;
  assign net_58386 = seg_14_15_local_g1_5_58386;
  assign net_58387 = seg_14_15_local_g1_6_58387;
  assign net_58391 = seg_14_15_local_g2_2_58391;
  assign net_58392 = seg_14_15_local_g2_3_58392;
  assign net_58395 = seg_14_15_local_g2_6_58395;
  assign net_58396 = seg_14_15_local_g2_7_58396;
  assign net_58397 = seg_14_15_local_g3_0_58397;
  assign net_58398 = seg_14_15_local_g3_1_58398;
  assign net_58402 = seg_14_15_local_g3_5_58402;
  assign net_58403 = seg_14_15_local_g3_6_58403;
  assign net_58404 = seg_14_15_local_g3_7_58404;
  assign net_58498 = seg_14_16_local_g0_2_58498;
  assign net_58500 = seg_14_16_local_g0_4_58500;
  assign net_58501 = seg_14_16_local_g0_5_58501;
  assign net_58504 = seg_14_16_local_g1_0_58504;
  assign net_58509 = seg_14_16_local_g1_5_58509;
  assign net_58511 = seg_14_16_local_g1_7_58511;
  assign net_58513 = seg_14_16_local_g2_1_58513;
  assign net_58517 = seg_14_16_local_g2_5_58517;
  assign net_58518 = seg_14_16_local_g2_6_58518;
  assign net_58520 = seg_14_16_local_g3_0_58520;
  assign net_58521 = seg_14_16_local_g3_1_58521;
  assign net_58523 = seg_14_16_local_g3_3_58523;
  assign net_58620 = seg_14_17_local_g0_1_58620;
  assign net_58630 = seg_14_17_local_g1_3_58630;
  assign net_58633 = seg_14_17_local_g1_6_58633;
  assign net_58644 = seg_14_17_local_g3_1_58644;
  assign net_58645 = seg_14_17_local_g3_2_58645;
  assign net_58650 = seg_14_17_local_g3_7_58650;
  assign net_58745 = seg_14_18_local_g0_3_58745;
  assign net_58747 = seg_14_18_local_g0_5_58747;
  assign net_58749 = seg_14_18_local_g0_7_58749;
  assign net_58753 = seg_14_18_local_g1_3_58753;
  assign net_58758 = seg_14_18_local_g2_0_58758;
  assign net_58759 = seg_14_18_local_g2_1_58759;
  assign net_58760 = seg_14_18_local_g2_2_58760;
  assign net_58761 = seg_14_18_local_g2_3_58761;
  assign net_58763 = seg_14_18_local_g2_5_58763;
  assign net_58764 = seg_14_18_local_g2_6_58764;
  assign net_58766 = seg_14_18_local_g3_0_58766;
  assign net_58767 = seg_14_18_local_g3_1_58767;
  assign net_58769 = seg_14_18_local_g3_3_58769;
  assign net_58865 = seg_14_19_local_g0_0_58865;
  assign net_58867 = seg_14_19_local_g0_2_58867;
  assign net_58873 = seg_14_19_local_g1_0_58873;
  assign net_58875 = seg_14_19_local_g1_2_58875;
  assign net_58877 = seg_14_19_local_g1_4_58877;
  assign net_58884 = seg_14_19_local_g2_3_58884;
  assign net_58892 = seg_14_19_local_g3_3_58892;
  assign net_58894 = seg_14_19_local_g3_5_58894;
  assign net_58988 = seg_14_20_local_g0_0_58988;
  assign net_58990 = seg_14_20_local_g0_2_58990;
  assign net_58991 = seg_14_20_local_g0_3_58991;
  assign net_58992 = seg_14_20_local_g0_4_58992;
  assign net_58993 = seg_14_20_local_g0_5_58993;
  assign net_58994 = seg_14_20_local_g0_6_58994;
  assign net_58995 = seg_14_20_local_g0_7_58995;
  assign net_58999 = seg_14_20_local_g1_3_58999;
  assign net_59002 = seg_14_20_local_g1_6_59002;
  assign net_59004 = seg_14_20_local_g2_0_59004;
  assign net_59005 = seg_14_20_local_g2_1_59005;
  assign net_59014 = seg_14_20_local_g3_2_59014;
  assign net_59016 = seg_14_20_local_g3_4_59016;
  assign net_59017 = seg_14_20_local_g3_5_59017;
  assign net_59140 = seg_14_21_local_g3_5_59140;
  assign net_59735 = seg_14_26_local_g1_1_59735;
  assign net_59737 = seg_14_26_local_g1_3_59737;
  assign net_59753 = seg_14_26_local_g3_3_59753;
  assign net_59851 = seg_14_27_local_g0_2_59851;
  assign net_59859 = seg_14_27_local_g1_2_59859;
  assign net_59862 = seg_14_27_local_g1_5_59862;
  assign net_59867 = seg_14_27_local_g2_2_59867;
  assign net_59869 = seg_14_27_local_g2_4_59869;
  assign net_59870 = seg_14_27_local_g2_5_59870;
  assign net_59875 = seg_14_27_local_g3_2_59875;
  assign net_59879 = seg_14_27_local_g3_6_59879;
  assign net_59984 = seg_14_28_local_g1_4_59984;
  assign net_59988 = seg_14_28_local_g2_0_59988;
  assign net_6 = seg_16_21_glb_netwk_1_6;
  assign net_60604 = seg_15_2_local_g0_0_60604;
  assign net_60606 = seg_15_2_local_g0_2_60606;
  assign net_60610 = seg_15_2_local_g0_6_60610;
  assign net_60611 = seg_15_2_local_g0_7_60611;
  assign net_60614 = seg_15_2_local_g1_2_60614;
  assign net_60615 = seg_15_2_local_g1_3_60615;
  assign net_60628 = seg_15_2_local_g3_0_60628;
  assign net_60729 = seg_15_3_local_g0_2_60729;
  assign net_60732 = seg_15_3_local_g0_5_60732;
  assign net_60735 = seg_15_3_local_g1_0_60735;
  assign net_60736 = seg_15_3_local_g1_1_60736;
  assign net_60738 = seg_15_3_local_g1_3_60738;
  assign net_60739 = seg_15_3_local_g1_4_60739;
  assign net_60740 = seg_15_3_local_g1_5_60740;
  assign net_60747 = seg_15_3_local_g2_4_60747;
  assign net_60749 = seg_15_3_local_g2_6_60749;
  assign net_60753 = seg_15_3_local_g3_2_60753;
  assign net_60754 = seg_15_3_local_g3_3_60754;
  assign net_60758 = seg_15_3_local_g3_7_60758;
  assign net_61119 = seg_15_6_local_g2_7_61119;
  assign net_61123 = seg_15_6_local_g3_3_61123;
  assign net_61350 = seg_15_8_local_g1_0_61350;
  assign net_61353 = seg_15_8_local_g1_3_61353;
  assign net_61473 = seg_15_9_local_g1_0_61473;
  assign net_61476 = seg_15_9_local_g1_3_61476;
  assign net_61483 = seg_15_9_local_g2_2_61483;
  assign net_61485 = seg_15_9_local_g2_4_61485;
  assign net_61486 = seg_15_9_local_g2_5_61486;
  assign net_61588 = seg_15_10_local_g0_0_61588;
  assign net_61591 = seg_15_10_local_g0_3_61591;
  assign net_61592 = seg_15_10_local_g0_4_61592;
  assign net_61594 = seg_15_10_local_g0_6_61594;
  assign net_61596 = seg_15_10_local_g1_0_61596;
  assign net_61598 = seg_15_10_local_g1_2_61598;
  assign net_61599 = seg_15_10_local_g1_3_61599;
  assign net_61600 = seg_15_10_local_g1_4_61600;
  assign net_61601 = seg_15_10_local_g1_5_61601;
  assign net_61602 = seg_15_10_local_g1_6_61602;
  assign net_61609 = seg_15_10_local_g2_5_61609;
  assign net_61610 = seg_15_10_local_g2_6_61610;
  assign net_61613 = seg_15_10_local_g3_1_61613;
  assign net_61616 = seg_15_10_local_g3_4_61616;
  assign net_61617 = seg_15_10_local_g3_5_61617;
  assign net_61715 = seg_15_11_local_g0_4_61715;
  assign net_61716 = seg_15_11_local_g0_5_61716;
  assign net_61717 = seg_15_11_local_g0_6_61717;
  assign net_61719 = seg_15_11_local_g1_0_61719;
  assign net_61724 = seg_15_11_local_g1_5_61724;
  assign net_61726 = seg_15_11_local_g1_7_61726;
  assign net_61728 = seg_15_11_local_g2_1_61728;
  assign net_61729 = seg_15_11_local_g2_2_61729;
  assign net_61730 = seg_15_11_local_g2_3_61730;
  assign net_61731 = seg_15_11_local_g2_4_61731;
  assign net_61735 = seg_15_11_local_g3_0_61735;
  assign net_61736 = seg_15_11_local_g3_1_61736;
  assign net_61737 = seg_15_11_local_g3_2_61737;
  assign net_61738 = seg_15_11_local_g3_3_61738;
  assign net_61739 = seg_15_11_local_g3_4_61739;
  assign net_61740 = seg_15_11_local_g3_5_61740;
  assign net_61741 = seg_15_11_local_g3_6_61741;
  assign net_61837 = seg_15_12_local_g0_3_61837;
  assign net_61838 = seg_15_12_local_g0_4_61838;
  assign net_61841 = seg_15_12_local_g0_7_61841;
  assign net_61842 = seg_15_12_local_g1_0_61842;
  assign net_61845 = seg_15_12_local_g1_3_61845;
  assign net_61850 = seg_15_12_local_g2_0_61850;
  assign net_61851 = seg_15_12_local_g2_1_61851;
  assign net_61852 = seg_15_12_local_g2_2_61852;
  assign net_61854 = seg_15_12_local_g2_4_61854;
  assign net_61855 = seg_15_12_local_g2_5_61855;
  assign net_61856 = seg_15_12_local_g2_6_61856;
  assign net_61857 = seg_15_12_local_g2_7_61857;
  assign net_61860 = seg_15_12_local_g3_2_61860;
  assign net_61861 = seg_15_12_local_g3_3_61861;
  assign net_61862 = seg_15_12_local_g3_4_61862;
  assign net_61863 = seg_15_12_local_g3_5_61863;
  assign net_61864 = seg_15_12_local_g3_6_61864;
  assign net_61957 = seg_15_13_local_g0_0_61957;
  assign net_61961 = seg_15_13_local_g0_4_61961;
  assign net_61962 = seg_15_13_local_g0_5_61962;
  assign net_61963 = seg_15_13_local_g0_6_61963;
  assign net_61965 = seg_15_13_local_g1_0_61965;
  assign net_61966 = seg_15_13_local_g1_1_61966;
  assign net_61967 = seg_15_13_local_g1_2_61967;
  assign net_61968 = seg_15_13_local_g1_3_61968;
  assign net_61969 = seg_15_13_local_g1_4_61969;
  assign net_61970 = seg_15_13_local_g1_5_61970;
  assign net_61972 = seg_15_13_local_g1_7_61972;
  assign net_61973 = seg_15_13_local_g2_0_61973;
  assign net_61974 = seg_15_13_local_g2_1_61974;
  assign net_61976 = seg_15_13_local_g2_3_61976;
  assign net_61977 = seg_15_13_local_g2_4_61977;
  assign net_61978 = seg_15_13_local_g2_5_61978;
  assign net_61983 = seg_15_13_local_g3_2_61983;
  assign net_61984 = seg_15_13_local_g3_3_61984;
  assign net_61985 = seg_15_13_local_g3_4_61985;
  assign net_61986 = seg_15_13_local_g3_5_61986;
  assign net_62081 = seg_15_14_local_g0_1_62081;
  assign net_62082 = seg_15_14_local_g0_2_62082;
  assign net_62083 = seg_15_14_local_g0_3_62083;
  assign net_62086 = seg_15_14_local_g0_6_62086;
  assign net_62089 = seg_15_14_local_g1_1_62089;
  assign net_62090 = seg_15_14_local_g1_2_62090;
  assign net_62092 = seg_15_14_local_g1_4_62092;
  assign net_62094 = seg_15_14_local_g1_6_62094;
  assign net_62095 = seg_15_14_local_g1_7_62095;
  assign net_62096 = seg_15_14_local_g2_0_62096;
  assign net_62098 = seg_15_14_local_g2_2_62098;
  assign net_62100 = seg_15_14_local_g2_4_62100;
  assign net_62101 = seg_15_14_local_g2_5_62101;
  assign net_62105 = seg_15_14_local_g3_1_62105;
  assign net_62111 = seg_15_14_local_g3_7_62111;
  assign net_62204 = seg_15_15_local_g0_1_62204;
  assign net_62206 = seg_15_15_local_g0_3_62206;
  assign net_62208 = seg_15_15_local_g0_5_62208;
  assign net_62209 = seg_15_15_local_g0_6_62209;
  assign net_62210 = seg_15_15_local_g0_7_62210;
  assign net_62217 = seg_15_15_local_g1_6_62217;
  assign net_62218 = seg_15_15_local_g1_7_62218;
  assign net_62220 = seg_15_15_local_g2_1_62220;
  assign net_62221 = seg_15_15_local_g2_2_62221;
  assign net_62224 = seg_15_15_local_g2_5_62224;
  assign net_62227 = seg_15_15_local_g3_0_62227;
  assign net_62229 = seg_15_15_local_g3_2_62229;
  assign net_62230 = seg_15_15_local_g3_3_62230;
  assign net_62232 = seg_15_15_local_g3_5_62232;
  assign net_62327 = seg_15_16_local_g0_1_62327;
  assign net_62331 = seg_15_16_local_g0_5_62331;
  assign net_62334 = seg_15_16_local_g1_0_62334;
  assign net_62337 = seg_15_16_local_g1_3_62337;
  assign net_62339 = seg_15_16_local_g1_5_62339;
  assign net_62340 = seg_15_16_local_g1_6_62340;
  assign net_62344 = seg_15_16_local_g2_2_62344;
  assign net_62346 = seg_15_16_local_g2_4_62346;
  assign net_62348 = seg_15_16_local_g2_6_62348;
  assign net_62350 = seg_15_16_local_g3_0_62350;
  assign net_62353 = seg_15_16_local_g3_3_62353;
  assign net_62354 = seg_15_16_local_g3_4_62354;
  assign net_62356 = seg_15_16_local_g3_6_62356;
  assign net_62456 = seg_15_17_local_g0_7_62456;
  assign net_62457 = seg_15_17_local_g1_0_62457;
  assign net_62458 = seg_15_17_local_g1_1_62458;
  assign net_62460 = seg_15_17_local_g1_3_62460;
  assign net_62467 = seg_15_17_local_g2_2_62467;
  assign net_62469 = seg_15_17_local_g2_4_62469;
  assign net_62470 = seg_15_17_local_g2_5_62470;
  assign net_62471 = seg_15_17_local_g2_6_62471;
  assign net_62472 = seg_15_17_local_g2_7_62472;
  assign net_62478 = seg_15_17_local_g3_5_62478;
  assign net_62479 = seg_15_17_local_g3_6_62479;
  assign net_62572 = seg_15_18_local_g0_0_62572;
  assign net_62573 = seg_15_18_local_g0_1_62573;
  assign net_62574 = seg_15_18_local_g0_2_62574;
  assign net_62578 = seg_15_18_local_g0_6_62578;
  assign net_62579 = seg_15_18_local_g0_7_62579;
  assign net_62582 = seg_15_18_local_g1_2_62582;
  assign net_62584 = seg_15_18_local_g1_4_62584;
  assign net_62588 = seg_15_18_local_g2_0_62588;
  assign net_62589 = seg_15_18_local_g2_1_62589;
  assign net_62592 = seg_15_18_local_g2_4_62592;
  assign net_62593 = seg_15_18_local_g2_5_62593;
  assign net_62597 = seg_15_18_local_g3_1_62597;
  assign net_62599 = seg_15_18_local_g3_3_62599;
  assign net_62600 = seg_15_18_local_g3_4_62600;
  assign net_62702 = seg_15_19_local_g0_7_62702;
  assign net_62703 = seg_15_19_local_g1_0_62703;
  assign net_62706 = seg_15_19_local_g1_3_62706;
  assign net_62715 = seg_15_19_local_g2_4_62715;
  assign net_62720 = seg_15_19_local_g3_1_62720;
  assign net_62722 = seg_15_19_local_g3_3_62722;
  assign net_62723 = seg_15_19_local_g3_4_62723;
  assign net_62724 = seg_15_19_local_g3_5_62724;
  assign net_62818 = seg_15_20_local_g0_0_62818;
  assign net_62821 = seg_15_20_local_g0_3_62821;
  assign net_62828 = seg_15_20_local_g1_2_62828;
  assign net_62829 = seg_15_20_local_g1_3_62829;
  assign net_62833 = seg_15_20_local_g1_7_62833;
  assign net_62834 = seg_15_20_local_g2_0_62834;
  assign net_62838 = seg_15_20_local_g2_4_62838;
  assign net_62844 = seg_15_20_local_g3_2_62844;
  assign net_62849 = seg_15_20_local_g3_7_62849;
  assign net_62956 = seg_15_21_local_g1_7_62956;
  assign net_62967 = seg_15_21_local_g3_2_62967;
  assign net_63068 = seg_15_22_local_g0_4_63068;
  assign net_63079 = seg_15_22_local_g1_7_63079;
  assign net_63091 = seg_15_22_local_g3_3_63091;
  assign net_63191 = seg_15_23_local_g0_4_63191;
  assign net_63192 = seg_15_23_local_g0_5_63192;
  assign net_63200 = seg_15_23_local_g1_5_63200;
  assign net_63204 = seg_15_23_local_g2_1_63204;
  assign net_63205 = seg_15_23_local_g2_2_63205;
  assign net_63439 = seg_15_25_local_g0_6_63439;
  assign net_63444 = seg_15_25_local_g1_3_63444;
  assign net_63683 = seg_15_27_local_g0_4_63683;
  assign net_63710 = seg_15_27_local_g3_7_63710;
  assign net_63807 = seg_15_28_local_g0_5_63807;
  assign net_63819 = seg_15_28_local_g2_1_63819;
  assign net_63823 = seg_15_28_local_g2_5_63823;
  assign net_63824 = seg_15_28_local_g2_6_63824;
  assign net_63829 = seg_15_28_local_g3_3_63829;
  assign net_63830 = seg_15_28_local_g3_4_63830;
  assign net_63831 = seg_15_28_local_g3_5_63831;
  assign net_63928 = seg_15_29_local_g0_3_63928;
  assign net_63930 = seg_15_29_local_g0_5_63930;
  assign net_63934 = seg_15_29_local_g1_1_63934;
  assign net_63936 = seg_15_29_local_g1_3_63936;
  assign net_63938 = seg_15_29_local_g1_5_63938;
  assign net_63939 = seg_15_29_local_g1_6_63939;
  assign net_63954 = seg_15_29_local_g3_5_63954;
  assign net_64436 = seg_16_2_local_g0_1_64436;
  assign net_64443 = seg_16_2_local_g1_0_64443;
  assign net_64444 = seg_16_2_local_g1_1_64444;
  assign net_64449 = seg_16_2_local_g1_6_64449;
  assign net_64455 = seg_16_2_local_g2_4_64455;
  assign net_64458 = seg_16_2_local_g2_7_64458;
  assign net_64461 = seg_16_2_local_g3_2_64461;
  assign net_64462 = seg_16_2_local_g3_3_64462;
  assign net_64466 = seg_16_2_local_g3_7_64466;
  assign net_64814 = seg_16_5_local_g1_2_64814;
  assign net_64818 = seg_16_5_local_g1_6_64818;
  assign net_64820 = seg_16_5_local_g2_0_64820;
  assign net_64827 = seg_16_5_local_g2_7_64827;
  assign net_64829 = seg_16_5_local_g3_1_64829;
  assign net_64830 = seg_16_5_local_g3_2_64830;
  assign net_64831 = seg_16_5_local_g3_3_64831;
  assign net_64834 = seg_16_5_local_g3_6_64834;
  assign net_64943 = seg_16_6_local_g2_0_64943;
  assign net_65298 = seg_16_9_local_g0_2_65298;
  assign net_65302 = seg_16_9_local_g0_6_65302;
  assign net_65304 = seg_16_9_local_g1_0_65304;
  assign net_65307 = seg_16_9_local_g1_3_65307;
  assign net_65308 = seg_16_9_local_g1_4_65308;
  assign net_65315 = seg_16_9_local_g2_3_65315;
  assign net_65318 = seg_16_9_local_g2_6_65318;
  assign net_65321 = seg_16_9_local_g3_1_65321;
  assign net_65428 = seg_16_10_local_g1_1_65428;
  assign net_65547 = seg_16_11_local_g0_5_65547;
  assign net_65548 = seg_16_11_local_g0_6_65548;
  assign net_65552 = seg_16_11_local_g1_2_65552;
  assign net_65566 = seg_16_11_local_g3_0_65566;
  assign net_65667 = seg_16_12_local_g0_2_65667;
  assign net_65674 = seg_16_12_local_g1_1_65674;
  assign net_65675 = seg_16_12_local_g1_2_65675;
  assign net_65677 = seg_16_12_local_g1_4_65677;
  assign net_65678 = seg_16_12_local_g1_5_65678;
  assign net_65679 = seg_16_12_local_g1_6_65679;
  assign net_65680 = seg_16_12_local_g1_7_65680;
  assign net_65683 = seg_16_12_local_g2_2_65683;
  assign net_65684 = seg_16_12_local_g2_3_65684;
  assign net_65686 = seg_16_12_local_g2_5_65686;
  assign net_65687 = seg_16_12_local_g2_6_65687;
  assign net_65688 = seg_16_12_local_g2_7_65688;
  assign net_65689 = seg_16_12_local_g3_0_65689;
  assign net_65693 = seg_16_12_local_g3_4_65693;
  assign net_65695 = seg_16_12_local_g3_6_65695;
  assign net_65790 = seg_16_13_local_g0_2_65790;
  assign net_65791 = seg_16_13_local_g0_3_65791;
  assign net_65792 = seg_16_13_local_g0_4_65792;
  assign net_65801 = seg_16_13_local_g1_5_65801;
  assign net_65806 = seg_16_13_local_g2_2_65806;
  assign net_65807 = seg_16_13_local_g2_3_65807;
  assign net_65812 = seg_16_13_local_g3_0_65812;
  assign net_65814 = seg_16_13_local_g3_2_65814;
  assign net_65917 = seg_16_14_local_g0_6_65917;
  assign net_65918 = seg_16_14_local_g0_7_65918;
  assign net_65935 = seg_16_14_local_g3_0_65935;
  assign net_65937 = seg_16_14_local_g3_2_65937;
  assign net_65942 = seg_16_14_local_g3_7_65942;
  assign net_66034 = seg_16_15_local_g0_0_66034;
  assign net_66035 = seg_16_15_local_g0_1_66035;
  assign net_66036 = seg_16_15_local_g0_2_66036;
  assign net_66040 = seg_16_15_local_g0_6_66040;
  assign net_66041 = seg_16_15_local_g0_7_66041;
  assign net_66042 = seg_16_15_local_g1_0_66042;
  assign net_66049 = seg_16_15_local_g1_7_66049;
  assign net_66050 = seg_16_15_local_g2_0_66050;
  assign net_66054 = seg_16_15_local_g2_4_66054;
  assign net_66055 = seg_16_15_local_g2_5_66055;
  assign net_66056 = seg_16_15_local_g2_6_66056;
  assign net_66057 = seg_16_15_local_g2_7_66057;
  assign net_66061 = seg_16_15_local_g3_3_66061;
  assign net_66062 = seg_16_15_local_g3_4_66062;
  assign net_66065 = seg_16_15_local_g3_7_66065;
  assign net_66158 = seg_16_16_local_g0_1_66158;
  assign net_66178 = seg_16_16_local_g2_5_66178;
  assign net_66181 = seg_16_16_local_g3_0_66181;
  assign net_66184 = seg_16_16_local_g3_3_66184;
  assign net_66281 = seg_16_17_local_g0_1_66281;
  assign net_66405 = seg_16_18_local_g0_2_66405;
  assign net_66408 = seg_16_18_local_g0_5_66408;
  assign net_66414 = seg_16_18_local_g1_3_66414;
  assign net_66415 = seg_16_18_local_g1_4_66415;
  assign net_66416 = seg_16_18_local_g1_5_66416;
  assign net_66422 = seg_16_18_local_g2_3_66422;
  assign net_66430 = seg_16_18_local_g3_3_66430;
  assign net_66433 = seg_16_18_local_g3_6_66433;
  assign net_66527 = seg_16_19_local_g0_1_66527;
  assign net_66528 = seg_16_19_local_g0_2_66528;
  assign net_66531 = seg_16_19_local_g0_5_66531;
  assign net_66533 = seg_16_19_local_g0_7_66533;
  assign net_66537 = seg_16_19_local_g1_3_66537;
  assign net_66538 = seg_16_19_local_g1_4_66538;
  assign net_66543 = seg_16_19_local_g2_1_66543;
  assign net_66546 = seg_16_19_local_g2_4_66546;
  assign net_66553 = seg_16_19_local_g3_3_66553;
  assign net_66554 = seg_16_19_local_g3_4_66554;
  assign net_66557 = seg_16_19_local_g3_7_66557;
  assign net_66650 = seg_16_20_local_g0_1_66650;
  assign net_66652 = seg_16_20_local_g0_3_66652;
  assign net_66653 = seg_16_20_local_g0_4_66653;
  assign net_66656 = seg_16_20_local_g0_7_66656;
  assign net_66658 = seg_16_20_local_g1_1_66658;
  assign net_66660 = seg_16_20_local_g1_3_66660;
  assign net_66661 = seg_16_20_local_g1_4_66661;
  assign net_66664 = seg_16_20_local_g1_7_66664;
  assign net_66667 = seg_16_20_local_g2_2_66667;
  assign net_66674 = seg_16_20_local_g3_1_66674;
  assign net_66675 = seg_16_20_local_g3_2_66675;
  assign net_66676 = seg_16_20_local_g3_3_66676;
  assign net_66797 = seg_16_21_local_g3_1_66797;
  assign net_67633 = seg_16_28_local_g0_0_67633;
  assign net_67635 = seg_16_28_local_g0_2_67635;
  assign net_67637 = seg_16_28_local_g0_4_67637;
  assign net_67642 = seg_16_28_local_g1_1_67642;
  assign net_67643 = seg_16_28_local_g1_2_67643;
  assign net_67645 = seg_16_28_local_g1_4_67645;
  assign net_67647 = seg_16_28_local_g1_6_67647;
  assign net_67649 = seg_16_28_local_g2_0_67649;
  assign net_67650 = seg_16_28_local_g2_1_67650;
  assign net_67654 = seg_16_28_local_g2_5_67654;
  assign net_67656 = seg_16_28_local_g2_7_67656;
  assign net_67657 = seg_16_28_local_g3_0_67657;
  assign net_67660 = seg_16_28_local_g3_3_67660;
  assign net_67757 = seg_16_29_local_g0_1_67757;
  assign net_67758 = seg_16_29_local_g0_2_67758;
  assign net_67759 = seg_16_29_local_g0_3_67759;
  assign net_67761 = seg_16_29_local_g0_5_67761;
  assign net_67765 = seg_16_29_local_g1_1_67765;
  assign net_67767 = seg_16_29_local_g1_3_67767;
  assign net_67770 = seg_16_29_local_g1_6_67770;
  assign net_67772 = seg_16_29_local_g2_0_67772;
  assign net_67774 = seg_16_29_local_g2_2_67774;
  assign net_67778 = seg_16_29_local_g2_6_67778;
  assign net_68056 = seg_17_0_local_g1_3_68056;
  assign net_68058 = seg_17_0_local_g1_5_68058;
  assign net_68638 = seg_17_5_local_g0_3_68638;
  assign net_68645 = seg_17_5_local_g1_2_68645;
  assign net_68646 = seg_17_5_local_g1_3_68646;
  assign net_68647 = seg_17_5_local_g1_4_68647;
  assign net_68648 = seg_17_5_local_g1_5_68648;
  assign net_68649 = seg_17_5_local_g1_6_68649;
  assign net_68650 = seg_17_5_local_g1_7_68650;
  assign net_68651 = seg_17_5_local_g2_0_68651;
  assign net_68655 = seg_17_5_local_g2_4_68655;
  assign net_68659 = seg_17_5_local_g3_0_68659;
  assign net_68662 = seg_17_5_local_g3_3_68662;
  assign net_68666 = seg_17_5_local_g3_7_68666;
  assign net_68758 = seg_17_6_local_g0_0_68758;
  assign net_68759 = seg_17_6_local_g0_1_68759;
  assign net_68764 = seg_17_6_local_g0_6_68764;
  assign net_68766 = seg_17_6_local_g1_0_68766;
  assign net_68768 = seg_17_6_local_g1_2_68768;
  assign net_68769 = seg_17_6_local_g1_3_68769;
  assign net_68771 = seg_17_6_local_g1_5_68771;
  assign net_68773 = seg_17_6_local_g1_7_68773;
  assign net_68774 = seg_17_6_local_g2_0_68774;
  assign net_68781 = seg_17_6_local_g2_7_68781;
  assign net_68782 = seg_17_6_local_g3_0_68782;
  assign net_68787 = seg_17_6_local_g3_5_68787;
  assign net_69151 = seg_17_9_local_g3_0_69151;
  assign net_69503 = seg_17_12_local_g0_7_69503;
  assign net_69525 = seg_17_12_local_g3_5_69525;
  assign net_69619 = seg_17_13_local_g0_0_69619;
  assign net_69623 = seg_17_13_local_g0_4_69623;
  assign net_69627 = seg_17_13_local_g1_0_69627;
  assign net_69629 = seg_17_13_local_g1_2_69629;
  assign net_69630 = seg_17_13_local_g1_3_69630;
  assign net_69742 = seg_17_14_local_g0_0_69742;
  assign net_69747 = seg_17_14_local_g0_5_69747;
  assign net_69749 = seg_17_14_local_g0_7_69749;
  assign net_69750 = seg_17_14_local_g1_0_69750;
  assign net_69753 = seg_17_14_local_g1_3_69753;
  assign net_69754 = seg_17_14_local_g1_4_69754;
  assign net_69756 = seg_17_14_local_g1_6_69756;
  assign net_69760 = seg_17_14_local_g2_2_69760;
  assign net_69763 = seg_17_14_local_g2_5_69763;
  assign net_69865 = seg_17_15_local_g0_0_69865;
  assign net_69867 = seg_17_15_local_g0_2_69867;
  assign net_69873 = seg_17_15_local_g1_0_69873;
  assign net_69875 = seg_17_15_local_g1_2_69875;
  assign net_69877 = seg_17_15_local_g1_4_69877;
  assign net_69878 = seg_17_15_local_g1_5_69878;
  assign net_69879 = seg_17_15_local_g1_6_69879;
  assign net_69880 = seg_17_15_local_g1_7_69880;
  assign net_70003 = seg_17_16_local_g1_7_70003;
  assign net_70014 = seg_17_16_local_g3_2_70014;
  assign net_70017 = seg_17_16_local_g3_5_70017;
  assign net_70112 = seg_17_17_local_g0_1_70112;
  assign net_70113 = seg_17_17_local_g0_2_70113;
  assign net_70120 = seg_17_17_local_g1_1_70120;
  assign net_70121 = seg_17_17_local_g1_2_70121;
  assign net_70123 = seg_17_17_local_g1_4_70123;
  assign net_70124 = seg_17_17_local_g1_5_70124;
  assign net_70128 = seg_17_17_local_g2_1_70128;
  assign net_70136 = seg_17_17_local_g3_1_70136;
  assign net_70137 = seg_17_17_local_g3_2_70137;
  assign net_70138 = seg_17_17_local_g3_3_70138;
  assign net_70140 = seg_17_17_local_g3_5_70140;
  assign net_70236 = seg_17_18_local_g0_2_70236;
  assign net_70239 = seg_17_18_local_g0_5_70239;
  assign net_70243 = seg_17_18_local_g1_1_70243;
  assign net_70245 = seg_17_18_local_g1_3_70245;
  assign net_70247 = seg_17_18_local_g1_5_70247;
  assign net_70248 = seg_17_18_local_g1_6_70248;
  assign net_70254 = seg_17_18_local_g2_4_70254;
  assign net_70358 = seg_17_19_local_g0_1_70358;
  assign net_70362 = seg_17_19_local_g0_5_70362;
  assign net_70363 = seg_17_19_local_g0_6_70363;
  assign net_70365 = seg_17_19_local_g1_0_70365;
  assign net_70371 = seg_17_19_local_g1_6_70371;
  assign net_70374 = seg_17_19_local_g2_1_70374;
  assign net_70375 = seg_17_19_local_g2_2_70375;
  assign net_70376 = seg_17_19_local_g2_3_70376;
  assign net_70379 = seg_17_19_local_g2_6_70379;
  assign net_70382 = seg_17_19_local_g3_1_70382;
  assign net_70385 = seg_17_19_local_g3_4_70385;
  assign net_70388 = seg_17_19_local_g3_7_70388;
  assign net_70489 = seg_17_20_local_g1_1_70489;
  assign net_70493 = seg_17_20_local_g1_5_70493;
  assign net_70494 = seg_17_20_local_g1_6_70494;
  assign net_70497 = seg_17_20_local_g2_1_70497;
  assign net_70501 = seg_17_20_local_g2_5_70501;
  assign net_70502 = seg_17_20_local_g2_6_70502;
  assign net_70503 = seg_17_20_local_g2_7_70503;
  assign net_70507 = seg_17_20_local_g3_3_70507;
  assign net_70508 = seg_17_20_local_g3_4_70508;
  assign net_70605 = seg_17_21_local_g0_2_70605;
  assign net_70606 = seg_17_21_local_g0_3_70606;
  assign net_70620 = seg_17_21_local_g2_1_70620;
  assign net_71604 = seg_17_29_local_g2_1_71604;
  assign net_71608 = seg_17_29_local_g2_5_71608;
  assign net_71609 = seg_17_29_local_g2_6_71609;
  assign net_71614 = seg_17_29_local_g3_3_71614;
  assign net_71851 = seg_17_31_local_g0_5_71851;
  assign net_71859 = seg_17_31_local_g1_5_71859;
  assign net_71878 = seg_18_0_local_g0_2_71878;
  assign net_71885 = seg_18_0_local_g1_1_71885;
  assign net_72466 = seg_18_5_local_g0_0_72466;
  assign net_72479 = seg_18_5_local_g1_5_72479;
  assign net_72484 = seg_18_5_local_g2_2_72484;
  assign net_72485 = seg_18_5_local_g2_3_72485;
  assign net_72495 = seg_18_5_local_g3_5_72495;
  assign net_72497 = seg_18_5_local_g3_7_72497;
  assign net_72593 = seg_18_6_local_g0_4_72593;
  assign net_72594 = seg_18_6_local_g0_5_72594;
  assign net_72596 = seg_18_6_local_g0_7_72596;
  assign net_72597 = seg_18_6_local_g1_0_72597;
  assign net_72600 = seg_18_6_local_g1_3_72600;
  assign net_72601 = seg_18_6_local_g1_4_72601;
  assign net_72602 = seg_18_6_local_g1_5_72602;
  assign net_72604 = seg_18_6_local_g1_7_72604;
  assign net_72605 = seg_18_6_local_g2_0_72605;
  assign net_72607 = seg_18_6_local_g2_2_72607;
  assign net_72610 = seg_18_6_local_g2_5_72610;
  assign net_72612 = seg_18_6_local_g2_7_72612;
  assign net_72613 = seg_18_6_local_g3_0_72613;
  assign net_72618 = seg_18_6_local_g3_5_72618;
  assign net_73084 = seg_18_10_local_g0_3_73084;
  assign net_73085 = seg_18_10_local_g0_4_73085;
  assign net_73090 = seg_18_10_local_g1_1_73090;
  assign net_73105 = seg_18_10_local_g3_0_73105;
  assign net_73330 = seg_18_12_local_g0_3_73330;
  assign net_73354 = seg_18_12_local_g3_3_73354;
  assign net_73355 = seg_18_12_local_g3_4_73355;
  assign net_73452 = seg_18_13_local_g0_2_73452;
  assign net_73453 = seg_18_13_local_g0_3_73453;
  assign net_73454 = seg_18_13_local_g0_4_73454;
  assign net_73461 = seg_18_13_local_g1_3_73461;
  assign net_73462 = seg_18_13_local_g1_4_73462;
  assign net_73467 = seg_18_13_local_g2_1_73467;
  assign net_73473 = seg_18_13_local_g2_7_73473;
  assign net_73475 = seg_18_13_local_g3_1_73475;
  assign net_73478 = seg_18_13_local_g3_4_73478;
  assign net_73479 = seg_18_13_local_g3_5_73479;
  assign net_73481 = seg_18_13_local_g3_7_73481;
  assign net_73574 = seg_18_14_local_g0_1_73574;
  assign net_73575 = seg_18_14_local_g0_2_73575;
  assign net_73576 = seg_18_14_local_g0_3_73576;
  assign net_73580 = seg_18_14_local_g0_7_73580;
  assign net_73582 = seg_18_14_local_g1_1_73582;
  assign net_73583 = seg_18_14_local_g1_2_73583;
  assign net_73585 = seg_18_14_local_g1_4_73585;
  assign net_73588 = seg_18_14_local_g1_7_73588;
  assign net_73589 = seg_18_14_local_g2_0_73589;
  assign net_73590 = seg_18_14_local_g2_1_73590;
  assign net_73591 = seg_18_14_local_g2_2_73591;
  assign net_73592 = seg_18_14_local_g2_3_73592;
  assign net_73595 = seg_18_14_local_g2_6_73595;
  assign net_73596 = seg_18_14_local_g2_7_73596;
  assign net_73599 = seg_18_14_local_g3_2_73599;
  assign net_73602 = seg_18_14_local_g3_5_73602;
  assign net_73604 = seg_18_14_local_g3_7_73604;
  assign net_73701 = seg_18_15_local_g0_5_73701;
  assign net_73713 = seg_18_15_local_g2_1_73713;
  assign net_73717 = seg_18_15_local_g2_5_73717;
  assign net_73722 = seg_18_15_local_g3_2_73722;
  assign net_73723 = seg_18_15_local_g3_3_73723;
  assign net_73724 = seg_18_15_local_g3_4_73724;
  assign net_73725 = seg_18_15_local_g3_5_73725;
  assign net_73845 = seg_18_16_local_g3_2_73845;
  assign net_73849 = seg_18_16_local_g3_6_73849;
  assign net_73946 = seg_18_17_local_g0_4_73946;
  assign net_73948 = seg_18_17_local_g0_6_73948;
  assign net_73950 = seg_18_17_local_g1_0_73950;
  assign net_73953 = seg_18_17_local_g1_3_73953;
  assign net_73955 = seg_18_17_local_g1_5_73955;
  assign net_73956 = seg_18_17_local_g1_6_73956;
  assign net_73962 = seg_18_17_local_g2_4_73962;
  assign net_73965 = seg_18_17_local_g2_7_73965;
  assign net_73969 = seg_18_17_local_g3_3_73969;
  assign net_73970 = seg_18_17_local_g3_4_73970;
  assign net_73971 = seg_18_17_local_g3_5_73971;
  assign net_74065 = seg_18_18_local_g0_0_74065;
  assign net_74068 = seg_18_18_local_g0_3_74068;
  assign net_74070 = seg_18_18_local_g0_5_74070;
  assign net_74072 = seg_18_18_local_g0_7_74072;
  assign net_74074 = seg_18_18_local_g1_1_74074;
  assign net_74076 = seg_18_18_local_g1_3_74076;
  assign net_74077 = seg_18_18_local_g1_4_74077;
  assign net_74080 = seg_18_18_local_g1_7_74080;
  assign net_74082 = seg_18_18_local_g2_1_74082;
  assign net_74083 = seg_18_18_local_g2_2_74083;
  assign net_74084 = seg_18_18_local_g2_3_74084;
  assign net_74086 = seg_18_18_local_g2_5_74086;
  assign net_74091 = seg_18_18_local_g3_2_74091;
  assign net_74092 = seg_18_18_local_g3_3_74092;
  assign net_74195 = seg_18_19_local_g0_7_74195;
  assign net_74320 = seg_18_20_local_g1_1_74320;
  assign net_75679 = seg_18_31_local_g0_2_75679;
  assign net_75682 = seg_18_31_local_g0_5_75682;
  assign net_77027 = seg_19_13_local_g0_0_77027;
  assign net_77030 = seg_19_13_local_g0_3_77030;
  assign net_77031 = seg_19_13_local_g0_4_77031;
  assign net_77033 = seg_19_13_local_g0_6_77033;
  assign net_77034 = seg_19_13_local_g0_7_77034;
  assign net_77035 = seg_19_13_local_g1_0_77035;
  assign net_77036 = seg_19_13_local_g1_1_77036;
  assign net_77038 = seg_19_13_local_g1_3_77038;
  assign net_77039 = seg_19_13_local_g1_4_77039;
  assign net_77040 = seg_19_13_local_g1_5_77040;
  assign net_77042 = seg_19_13_local_g1_7_77042;
  assign net_77044 = seg_19_13_local_g2_1_77044;
  assign net_77048 = seg_19_13_local_g2_5_77048;
  assign net_77049 = seg_19_13_local_g2_6_77049;
  assign net_77050 = seg_19_13_local_g2_7_77050;
  assign net_77054 = seg_19_13_local_g3_3_77054;
  assign net_77056 = seg_19_13_local_g3_5_77056;
  assign net_77057 = seg_19_13_local_g3_6_77057;
  assign net_77129 = seg_19_14_local_g0_0_77129;
  assign net_77130 = seg_19_14_local_g0_1_77130;
  assign net_77131 = seg_19_14_local_g0_2_77131;
  assign net_77132 = seg_19_14_local_g0_3_77132;
  assign net_77133 = seg_19_14_local_g0_4_77133;
  assign net_77134 = seg_19_14_local_g0_5_77134;
  assign net_77135 = seg_19_14_local_g0_6_77135;
  assign net_77137 = seg_19_14_local_g1_0_77137;
  assign net_77141 = seg_19_14_local_g1_4_77141;
  assign net_77142 = seg_19_14_local_g1_5_77142;
  assign net_77147 = seg_19_14_local_g2_2_77147;
  assign net_77150 = seg_19_14_local_g2_5_77150;
  assign net_77151 = seg_19_14_local_g2_6_77151;
  assign net_77152 = seg_19_14_local_g2_7_77152;
  assign net_77156 = seg_19_14_local_g3_3_77156;
  assign net_77157 = seg_19_14_local_g3_4_77157;
  assign net_77158 = seg_19_14_local_g3_5_77158;
  assign net_77160 = seg_19_14_local_g3_7_77160;
  assign net_77231 = seg_19_15_local_g0_0_77231;
  assign net_77232 = seg_19_15_local_g0_1_77232;
  assign net_77233 = seg_19_15_local_g0_2_77233;
  assign net_77234 = seg_19_15_local_g0_3_77234;
  assign net_77235 = seg_19_15_local_g0_4_77235;
  assign net_77236 = seg_19_15_local_g0_5_77236;
  assign net_77239 = seg_19_15_local_g1_0_77239;
  assign net_77240 = seg_19_15_local_g1_1_77240;
  assign net_77246 = seg_19_15_local_g1_7_77246;
  assign net_77247 = seg_19_15_local_g2_0_77247;
  assign net_77248 = seg_19_15_local_g2_1_77248;
  assign net_77251 = seg_19_15_local_g2_4_77251;
  assign net_77252 = seg_19_15_local_g2_5_77252;
  assign net_77254 = seg_19_15_local_g2_7_77254;
  assign net_77258 = seg_19_15_local_g3_3_77258;
  assign net_77260 = seg_19_15_local_g3_5_77260;
  assign net_77261 = seg_19_15_local_g3_6_77261;
  assign net_77262 = seg_19_15_local_g3_7_77262;
  assign net_77334 = seg_19_16_local_g0_1_77334;
  assign net_77339 = seg_19_16_local_g0_6_77339;
  assign net_77342 = seg_19_16_local_g1_1_77342;
  assign net_77343 = seg_19_16_local_g1_2_77343;
  assign net_77346 = seg_19_16_local_g1_5_77346;
  assign net_77349 = seg_19_16_local_g2_0_77349;
  assign net_77351 = seg_19_16_local_g2_2_77351;
  assign net_77353 = seg_19_16_local_g2_4_77353;
  assign net_77354 = seg_19_16_local_g2_5_77354;
  assign net_77356 = seg_19_16_local_g2_7_77356;
  assign net_77357 = seg_19_16_local_g3_0_77357;
  assign net_77358 = seg_19_16_local_g3_1_77358;
  assign net_77359 = seg_19_16_local_g3_2_77359;
  assign net_77360 = seg_19_16_local_g3_3_77360;
  assign net_77361 = seg_19_16_local_g3_4_77361;
  assign net_77362 = seg_19_16_local_g3_5_77362;
  assign net_77363 = seg_19_16_local_g3_6_77363;
  assign net_77364 = seg_19_16_local_g3_7_77364;
  assign net_77435 = seg_19_17_local_g0_0_77435;
  assign net_77436 = seg_19_17_local_g0_1_77436;
  assign net_77437 = seg_19_17_local_g0_2_77437;
  assign net_77439 = seg_19_17_local_g0_4_77439;
  assign net_77440 = seg_19_17_local_g0_5_77440;
  assign net_77446 = seg_19_17_local_g1_3_77446;
  assign net_77447 = seg_19_17_local_g1_4_77447;
  assign net_77449 = seg_19_17_local_g1_6_77449;
  assign net_77450 = seg_19_17_local_g1_7_77450;
  assign net_77452 = seg_19_17_local_g2_1_77452;
  assign net_77453 = seg_19_17_local_g2_2_77453;
  assign net_77456 = seg_19_17_local_g2_5_77456;
  assign net_77457 = seg_19_17_local_g2_6_77457;
  assign net_77461 = seg_19_17_local_g3_2_77461;
  assign net_77462 = seg_19_17_local_g3_3_77462;
  assign net_77464 = seg_19_17_local_g3_5_77464;
  assign net_77466 = seg_19_17_local_g3_7_77466;
  assign net_77538 = seg_19_18_local_g0_1_77538;
  assign net_77539 = seg_19_18_local_g0_2_77539;
  assign net_77541 = seg_19_18_local_g0_4_77541;
  assign net_77542 = seg_19_18_local_g0_5_77542;
  assign net_77545 = seg_19_18_local_g1_0_77545;
  assign net_77548 = seg_19_18_local_g1_3_77548;
  assign net_77549 = seg_19_18_local_g1_4_77549;
  assign net_77550 = seg_19_18_local_g1_5_77550;
  assign net_77553 = seg_19_18_local_g2_0_77553;
  assign net_77555 = seg_19_18_local_g2_2_77555;
  assign net_77558 = seg_19_18_local_g2_5_77558;
  assign net_77559 = seg_19_18_local_g2_6_77559;
  assign net_77561 = seg_19_18_local_g3_0_77561;
  assign net_77562 = seg_19_18_local_g3_1_77562;
  assign net_77563 = seg_19_18_local_g3_2_77563;
  assign net_77564 = seg_19_18_local_g3_3_77564;
  assign net_77565 = seg_19_18_local_g3_4_77565;
  assign net_77568 = seg_19_18_local_g3_7_77568;
  assign net_79622 = seg_20_6_local_g0_2_79622;
  assign net_79624 = seg_20_6_local_g0_4_79624;
  assign net_79628 = seg_20_6_local_g1_0_79628;
  assign net_79630 = seg_20_6_local_g1_2_79630;
  assign net_79635 = seg_20_6_local_g1_7_79635;
  assign net_79638 = seg_20_6_local_g2_2_79638;
  assign net_79641 = seg_20_6_local_g2_5_79641;
  assign net_79646 = seg_20_6_local_g3_2_79646;
  assign net_79649 = seg_20_6_local_g3_5_79649;
  assign net_79756 = seg_20_7_local_g1_5_79756;
  assign net_79761 = seg_20_7_local_g2_2_79761;
  assign net_79991 = seg_20_9_local_g0_2_79991;
  assign net_79997 = seg_20_9_local_g1_0_79997;
  assign net_8 = seg_17_20_glb_netwk_3_8;
  assign net_80000 = seg_20_9_local_g1_3_80000;
  assign net_80004 = seg_20_9_local_g1_7_80004;
  assign net_80014 = seg_20_9_local_g3_1_80014;
  assign net_80114 = seg_20_10_local_g0_2_80114;
  assign net_80117 = seg_20_10_local_g0_5_80117;
  assign net_80119 = seg_20_10_local_g0_7_80119;
  assign net_80121 = seg_20_10_local_g1_1_80121;
  assign net_80122 = seg_20_10_local_g1_2_80122;
  assign net_80123 = seg_20_10_local_g1_3_80123;
  assign net_80125 = seg_20_10_local_g1_5_80125;
  assign net_80129 = seg_20_10_local_g2_1_80129;
  assign net_80132 = seg_20_10_local_g2_4_80132;
  assign net_80136 = seg_20_10_local_g3_0_80136;
  assign net_80137 = seg_20_10_local_g3_1_80137;
  assign net_80139 = seg_20_10_local_g3_3_80139;
  assign net_80140 = seg_20_10_local_g3_4_80140;
  assign net_80242 = seg_20_11_local_g0_7_80242;
  assign net_80359 = seg_20_12_local_g0_1_80359;
  assign net_80360 = seg_20_12_local_g0_2_80360;
  assign net_80364 = seg_20_12_local_g0_6_80364;
  assign net_80368 = seg_20_12_local_g1_2_80368;
  assign net_80369 = seg_20_12_local_g1_3_80369;
  assign net_80371 = seg_20_12_local_g1_5_80371;
  assign net_80372 = seg_20_12_local_g1_6_80372;
  assign net_80373 = seg_20_12_local_g1_7_80373;
  assign net_80375 = seg_20_12_local_g2_1_80375;
  assign net_80376 = seg_20_12_local_g2_2_80376;
  assign net_80377 = seg_20_12_local_g2_3_80377;
  assign net_80378 = seg_20_12_local_g2_4_80378;
  assign net_80379 = seg_20_12_local_g2_5_80379;
  assign net_80380 = seg_20_12_local_g2_6_80380;
  assign net_80381 = seg_20_12_local_g2_7_80381;
  assign net_80385 = seg_20_12_local_g3_3_80385;
  assign net_80388 = seg_20_12_local_g3_6_80388;
  assign net_80389 = seg_20_12_local_g3_7_80389;
  assign net_80481 = seg_20_13_local_g0_0_80481;
  assign net_80482 = seg_20_13_local_g0_1_80482;
  assign net_80483 = seg_20_13_local_g0_2_80483;
  assign net_80485 = seg_20_13_local_g0_4_80485;
  assign net_80486 = seg_20_13_local_g0_5_80486;
  assign net_80489 = seg_20_13_local_g1_0_80489;
  assign net_80491 = seg_20_13_local_g1_2_80491;
  assign net_80492 = seg_20_13_local_g1_3_80492;
  assign net_80493 = seg_20_13_local_g1_4_80493;
  assign net_80494 = seg_20_13_local_g1_5_80494;
  assign net_80495 = seg_20_13_local_g1_6_80495;
  assign net_80499 = seg_20_13_local_g2_2_80499;
  assign net_80501 = seg_20_13_local_g2_4_80501;
  assign net_80502 = seg_20_13_local_g2_5_80502;
  assign net_80503 = seg_20_13_local_g2_6_80503;
  assign net_80507 = seg_20_13_local_g3_2_80507;
  assign net_80509 = seg_20_13_local_g3_4_80509;
  assign net_80510 = seg_20_13_local_g3_5_80510;
  assign net_80511 = seg_20_13_local_g3_6_80511;
  assign net_80604 = seg_20_14_local_g0_0_80604;
  assign net_80605 = seg_20_14_local_g0_1_80605;
  assign net_80609 = seg_20_14_local_g0_5_80609;
  assign net_80611 = seg_20_14_local_g0_7_80611;
  assign net_80612 = seg_20_14_local_g1_0_80612;
  assign net_80613 = seg_20_14_local_g1_1_80613;
  assign net_80618 = seg_20_14_local_g1_6_80618;
  assign net_80619 = seg_20_14_local_g1_7_80619;
  assign net_80620 = seg_20_14_local_g2_0_80620;
  assign net_80622 = seg_20_14_local_g2_2_80622;
  assign net_80623 = seg_20_14_local_g2_3_80623;
  assign net_80624 = seg_20_14_local_g2_4_80624;
  assign net_80626 = seg_20_14_local_g2_6_80626;
  assign net_80628 = seg_20_14_local_g3_0_80628;
  assign net_80631 = seg_20_14_local_g3_3_80631;
  assign net_80635 = seg_20_14_local_g3_7_80635;
  assign net_80727 = seg_20_15_local_g0_0_80727;
  assign net_80729 = seg_20_15_local_g0_2_80729;
  assign net_80731 = seg_20_15_local_g0_4_80731;
  assign net_80735 = seg_20_15_local_g1_0_80735;
  assign net_80736 = seg_20_15_local_g1_1_80736;
  assign net_80738 = seg_20_15_local_g1_3_80738;
  assign net_80739 = seg_20_15_local_g1_4_80739;
  assign net_80740 = seg_20_15_local_g1_5_80740;
  assign net_80741 = seg_20_15_local_g1_6_80741;
  assign net_80743 = seg_20_15_local_g2_0_80743;
  assign net_80744 = seg_20_15_local_g2_1_80744;
  assign net_80745 = seg_20_15_local_g2_2_80745;
  assign net_80747 = seg_20_15_local_g2_4_80747;
  assign net_80749 = seg_20_15_local_g2_6_80749;
  assign net_80751 = seg_20_15_local_g3_0_80751;
  assign net_80752 = seg_20_15_local_g3_1_80752;
  assign net_80753 = seg_20_15_local_g3_2_80753;
  assign net_80755 = seg_20_15_local_g3_4_80755;
  assign net_80757 = seg_20_15_local_g3_6_80757;
  assign net_80855 = seg_20_16_local_g0_5_80855;
  assign net_80859 = seg_20_16_local_g1_1_80859;
  assign net_80862 = seg_20_16_local_g1_4_80862;
  assign net_80864 = seg_20_16_local_g1_6_80864;
  assign net_80868 = seg_20_16_local_g2_2_80868;
  assign net_80870 = seg_20_16_local_g2_4_80870;
  assign net_80871 = seg_20_16_local_g2_5_80871;
  assign net_80877 = seg_20_16_local_g3_3_80877;
  assign net_80881 = seg_20_16_local_g3_7_80881;
  assign net_80975 = seg_20_17_local_g0_2_80975;
  assign net_80976 = seg_20_17_local_g0_3_80976;
  assign net_80977 = seg_20_17_local_g0_4_80977;
  assign net_80978 = seg_20_17_local_g0_5_80978;
  assign net_80979 = seg_20_17_local_g0_6_80979;
  assign net_80980 = seg_20_17_local_g0_7_80980;
  assign net_80984 = seg_20_17_local_g1_3_80984;
  assign net_80985 = seg_20_17_local_g1_4_80985;
  assign net_80986 = seg_20_17_local_g1_5_80986;
  assign net_80987 = seg_20_17_local_g1_6_80987;
  assign net_80989 = seg_20_17_local_g2_0_80989;
  assign net_80990 = seg_20_17_local_g2_1_80990;
  assign net_80991 = seg_20_17_local_g2_2_80991;
  assign net_80992 = seg_20_17_local_g2_3_80992;
  assign net_80993 = seg_20_17_local_g2_4_80993;
  assign net_80995 = seg_20_17_local_g2_6_80995;
  assign net_80996 = seg_20_17_local_g2_7_80996;
  assign net_80997 = seg_20_17_local_g3_0_80997;
  assign net_80998 = seg_20_17_local_g3_1_80998;
  assign net_81001 = seg_20_17_local_g3_4_81001;
  assign net_81002 = seg_20_17_local_g3_5_81002;
  assign net_81003 = seg_20_17_local_g3_6_81003;
  assign net_81098 = seg_20_18_local_g0_2_81098;
  assign net_81099 = seg_20_18_local_g0_3_81099;
  assign net_81102 = seg_20_18_local_g0_6_81102;
  assign net_81103 = seg_20_18_local_g0_7_81103;
  assign net_81105 = seg_20_18_local_g1_1_81105;
  assign net_81107 = seg_20_18_local_g1_3_81107;
  assign net_81110 = seg_20_18_local_g1_6_81110;
  assign net_81111 = seg_20_18_local_g1_7_81111;
  assign net_81112 = seg_20_18_local_g2_0_81112;
  assign net_81115 = seg_20_18_local_g2_3_81115;
  assign net_81119 = seg_20_18_local_g2_7_81119;
  assign net_81120 = seg_20_18_local_g3_0_81120;
  assign net_81125 = seg_20_18_local_g3_5_81125;
  assign net_81236 = seg_20_19_local_g2_1_81236;
  assign net_81240 = seg_20_19_local_g2_5_81240;
  assign net_83456 = seg_21_6_local_g0_5_83456;
  assign net_83460 = seg_21_6_local_g1_1_83460;
  assign net_83466 = seg_21_6_local_g1_7_83466;
  assign net_83822 = seg_21_9_local_g0_2_83822;
  assign net_83828 = seg_21_9_local_g1_0_83828;
  assign net_83833 = seg_21_9_local_g1_5_83833;
  assign net_83835 = seg_21_9_local_g1_7_83835;
  assign net_83843 = seg_21_9_local_g2_7_83843;
  assign net_83849 = seg_21_9_local_g3_5_83849;
  assign net_83943 = seg_21_10_local_g0_0_83943;
  assign net_83945 = seg_21_10_local_g0_2_83945;
  assign net_83946 = seg_21_10_local_g0_3_83946;
  assign net_83947 = seg_21_10_local_g0_4_83947;
  assign net_83956 = seg_21_10_local_g1_5_83956;
  assign net_83963 = seg_21_10_local_g2_4_83963;
  assign net_83964 = seg_21_10_local_g2_5_83964;
  assign net_83967 = seg_21_10_local_g3_0_83967;
  assign net_83972 = seg_21_10_local_g3_5_83972;
  assign net_84189 = seg_21_12_local_g0_0_84189;
  assign net_84196 = seg_21_12_local_g0_7_84196;
  assign net_84197 = seg_21_12_local_g1_0_84197;
  assign net_84202 = seg_21_12_local_g1_5_84202;
  assign net_84204 = seg_21_12_local_g1_7_84204;
  assign net_84217 = seg_21_12_local_g3_4_84217;
  assign net_84313 = seg_21_13_local_g0_1_84313;
  assign net_84314 = seg_21_13_local_g0_2_84314;
  assign net_84316 = seg_21_13_local_g0_4_84316;
  assign net_84319 = seg_21_13_local_g0_7_84319;
  assign net_84321 = seg_21_13_local_g1_1_84321;
  assign net_84322 = seg_21_13_local_g1_2_84322;
  assign net_84324 = seg_21_13_local_g1_4_84324;
  assign net_84325 = seg_21_13_local_g1_5_84325;
  assign net_84326 = seg_21_13_local_g1_6_84326;
  assign net_84327 = seg_21_13_local_g1_7_84327;
  assign net_84328 = seg_21_13_local_g2_0_84328;
  assign net_84333 = seg_21_13_local_g2_5_84333;
  assign net_84334 = seg_21_13_local_g2_6_84334;
  assign net_84335 = seg_21_13_local_g2_7_84335;
  assign net_84338 = seg_21_13_local_g3_2_84338;
  assign net_84341 = seg_21_13_local_g3_5_84341;
  assign net_84342 = seg_21_13_local_g3_6_84342;
  assign net_84343 = seg_21_13_local_g3_7_84343;
  assign net_84436 = seg_21_14_local_g0_1_84436;
  assign net_84437 = seg_21_14_local_g0_2_84437;
  assign net_84438 = seg_21_14_local_g0_3_84438;
  assign net_84439 = seg_21_14_local_g0_4_84439;
  assign net_84441 = seg_21_14_local_g0_6_84441;
  assign net_84442 = seg_21_14_local_g0_7_84442;
  assign net_84443 = seg_21_14_local_g1_0_84443;
  assign net_84444 = seg_21_14_local_g1_1_84444;
  assign net_84445 = seg_21_14_local_g1_2_84445;
  assign net_84446 = seg_21_14_local_g1_3_84446;
  assign net_84447 = seg_21_14_local_g1_4_84447;
  assign net_84448 = seg_21_14_local_g1_5_84448;
  assign net_84450 = seg_21_14_local_g1_7_84450;
  assign net_84452 = seg_21_14_local_g2_1_84452;
  assign net_84453 = seg_21_14_local_g2_2_84453;
  assign net_84454 = seg_21_14_local_g2_3_84454;
  assign net_84455 = seg_21_14_local_g2_4_84455;
  assign net_84456 = seg_21_14_local_g2_5_84456;
  assign net_84458 = seg_21_14_local_g2_7_84458;
  assign net_84459 = seg_21_14_local_g3_0_84459;
  assign net_84462 = seg_21_14_local_g3_3_84462;
  assign net_84463 = seg_21_14_local_g3_4_84463;
  assign net_84465 = seg_21_14_local_g3_6_84465;
  assign net_84466 = seg_21_14_local_g3_7_84466;
  assign net_84558 = seg_21_15_local_g0_0_84558;
  assign net_84560 = seg_21_15_local_g0_2_84560;
  assign net_84561 = seg_21_15_local_g0_3_84561;
  assign net_84562 = seg_21_15_local_g0_4_84562;
  assign net_84563 = seg_21_15_local_g0_5_84563;
  assign net_84564 = seg_21_15_local_g0_6_84564;
  assign net_84566 = seg_21_15_local_g1_0_84566;
  assign net_84567 = seg_21_15_local_g1_1_84567;
  assign net_84568 = seg_21_15_local_g1_2_84568;
  assign net_84569 = seg_21_15_local_g1_3_84569;
  assign net_84570 = seg_21_15_local_g1_4_84570;
  assign net_84571 = seg_21_15_local_g1_5_84571;
  assign net_84572 = seg_21_15_local_g1_6_84572;
  assign net_84573 = seg_21_15_local_g1_7_84573;
  assign net_84575 = seg_21_15_local_g2_1_84575;
  assign net_84578 = seg_21_15_local_g2_4_84578;
  assign net_84581 = seg_21_15_local_g2_7_84581;
  assign net_84582 = seg_21_15_local_g3_0_84582;
  assign net_84583 = seg_21_15_local_g3_1_84583;
  assign net_84584 = seg_21_15_local_g3_2_84584;
  assign net_84585 = seg_21_15_local_g3_3_84585;
  assign net_84586 = seg_21_15_local_g3_4_84586;
  assign net_84589 = seg_21_15_local_g3_7_84589;
  assign net_84682 = seg_21_16_local_g0_1_84682;
  assign net_84686 = seg_21_16_local_g0_5_84686;
  assign net_84694 = seg_21_16_local_g1_5_84694;
  assign net_84696 = seg_21_16_local_g1_7_84696;
  assign net_84698 = seg_21_16_local_g2_1_84698;
  assign net_84706 = seg_21_16_local_g3_1_84706;
  assign net_84711 = seg_21_16_local_g3_6_84711;
  assign net_84806 = seg_21_17_local_g0_2_84806;
  assign net_84808 = seg_21_17_local_g0_4_84808;
  assign net_84812 = seg_21_17_local_g1_0_84812;
  assign net_84813 = seg_21_17_local_g1_1_84813;
  assign net_84814 = seg_21_17_local_g1_2_84814;
  assign net_84815 = seg_21_17_local_g1_3_84815;
  assign net_84817 = seg_21_17_local_g1_5_84817;
  assign net_84821 = seg_21_17_local_g2_1_84821;
  assign net_84822 = seg_21_17_local_g2_2_84822;
  assign net_84824 = seg_21_17_local_g2_4_84824;
  assign net_84825 = seg_21_17_local_g2_5_84825;
  assign net_84826 = seg_21_17_local_g2_6_84826;
  assign net_84827 = seg_21_17_local_g2_7_84827;
  assign net_84829 = seg_21_17_local_g3_1_84829;
  assign net_84830 = seg_21_17_local_g3_2_84830;
  assign net_84831 = seg_21_17_local_g3_3_84831;
  assign net_84832 = seg_21_17_local_g3_4_84832;
  assign net_84833 = seg_21_17_local_g3_5_84833;
  assign net_84834 = seg_21_17_local_g3_6_84834;
  assign net_84835 = seg_21_17_local_g3_7_84835;
  assign net_84928 = seg_21_18_local_g0_1_84928;
  assign net_84929 = seg_21_18_local_g0_2_84929;
  assign net_84930 = seg_21_18_local_g0_3_84930;
  assign net_84931 = seg_21_18_local_g0_4_84931;
  assign net_84935 = seg_21_18_local_g1_0_84935;
  assign net_84936 = seg_21_18_local_g1_1_84936;
  assign net_84938 = seg_21_18_local_g1_3_84938;
  assign net_84939 = seg_21_18_local_g1_4_84939;
  assign net_84940 = seg_21_18_local_g1_5_84940;
  assign net_84941 = seg_21_18_local_g1_6_84941;
  assign net_84952 = seg_21_18_local_g3_1_84952;
  assign net_84953 = seg_21_18_local_g3_2_84953;
  assign net_84955 = seg_21_18_local_g3_4_84955;
  assign net_84957 = seg_21_18_local_g3_6_84957;
  assign net_85064 = seg_21_19_local_g1_6_85064;
  assign net_86579 = seg_22_0_local_g1_2_86579;
  assign net_87652 = seg_22_9_local_g0_1_87652;
  assign net_87655 = seg_22_9_local_g0_4_87655;
  assign net_87669 = seg_22_9_local_g2_2_87669;
  assign net_88152 = seg_22_13_local_g1_1_88152;
  assign net_88166 = seg_22_13_local_g2_7_88166;
  assign net_88270 = seg_22_14_local_g0_4_88270;
  assign net_88278 = seg_22_14_local_g1_4_88278;
  assign net_88279 = seg_22_14_local_g1_5_88279;
  assign net_88417 = seg_22_15_local_g3_4_88417;
  assign net_88419 = seg_22_15_local_g3_6_88419;
  assign net_88534 = seg_22_16_local_g2_6_88534;
  assign net_88539 = seg_22_16_local_g3_3_88539;
  assign net_88636 = seg_22_17_local_g0_1_88636;
  assign net_88638 = seg_22_17_local_g0_3_88638;
  assign net_88639 = seg_22_17_local_g0_4_88639;
  assign net_88640 = seg_22_17_local_g0_5_88640;
  assign net_88642 = seg_22_17_local_g0_7_88642;
  assign net_88646 = seg_22_17_local_g1_3_88646;
  assign net_88647 = seg_22_17_local_g1_4_88647;
  assign net_88650 = seg_22_17_local_g1_7_88650;
  assign net_88656 = seg_22_17_local_g2_5_88656;
  assign net_91484 = seg_23_9_local_g0_2_91484;
  assign net_91491 = seg_23_9_local_g1_1_91491;
  assign net_91493 = seg_23_9_local_g1_3_91493;
  assign net_91495 = seg_23_9_local_g1_5_91495;
  assign net_91506 = seg_23_9_local_g3_0_91506;
  assign seg_10_10_lutff_2_out_38565 = net_38565;
  assign seg_10_10_neigh_op_lft_1_34733 = seg_9_10_lutff_1_out_34733;
  assign seg_10_10_sp4_h_l_43_27633 = seg_8_10_sp4_h_r_30_27633;
  assign seg_10_10_sp4_h_r_36_31037 = net_31037;
  assign seg_10_10_sp4_h_r_4_42535 = net_42535;
  assign seg_10_11_lutff_0_out_38686 = net_38686;
  assign seg_10_11_lutff_1_out_38687 = net_38687;
  assign seg_10_11_lutff_4_out_38690 = net_38690;
  assign seg_10_11_neigh_op_bnl_4_34736 = seg_9_10_lutff_4_out_34736;
  assign seg_10_11_neigh_op_bot_2_38565 = seg_10_10_lutff_2_out_38565;
  assign seg_10_11_neigh_op_lft_5_34860 = seg_9_11_lutff_5_out_34860;
  assign seg_10_11_neigh_op_rgt_2_42519 = seg_11_11_lutff_2_out_42519;
  assign seg_10_11_neigh_op_rgt_7_42524 = seg_11_11_lutff_7_out_42524;
  assign seg_10_11_sp4_r_v_b_37_42665 = net_42665;
  assign seg_10_12_lutff_1_out_38810 = net_38810;
  assign seg_10_12_lutff_5_out_38814 = net_38814;
  assign seg_10_12_lutff_7_out_38816 = net_38816;
  assign seg_10_12_neigh_op_bot_0_38686 = seg_10_11_lutff_0_out_38686;
  assign seg_10_12_neigh_op_bot_1_38687 = seg_10_11_lutff_1_out_38687;
  assign seg_10_12_neigh_op_bot_4_38690 = seg_10_11_lutff_4_out_38690;
  assign seg_10_12_neigh_op_rgt_6_42646 = seg_11_12_lutff_6_out_42646;
  assign seg_10_12_sp4_h_r_11_42778 = seg_13_12_sp4_h_r_46_42778;
  assign seg_10_12_sp4_h_r_12_38945 = net_38945;
  assign seg_10_12_sp4_h_r_4_42781 = net_42781;
  assign seg_10_12_sp4_h_r_6_42783 = net_42783;
  assign seg_10_12_sp4_h_r_8_42785 = net_42785;
  assign seg_10_12_sp4_r_v_b_35_42674 = seg_10_14_sp4_r_v_b_11_42674;
  assign seg_10_12_sp4_v_b_17_38715 = seg_9_10_sp4_r_v_b_41_38715;
  assign seg_10_12_sp4_v_b_45_38965 = seg_10_15_sp4_v_b_8_38965;
  assign seg_10_13_lutff_1_out_38933 = net_38933;
  assign seg_10_13_lutff_2_out_38934 = net_38934;
  assign seg_10_13_lutff_4_out_38936 = net_38936;
  assign seg_10_13_lutff_5_out_38937 = net_38937;
  assign seg_10_13_lutff_6_out_38938 = net_38938;
  assign seg_10_13_lutff_7_out_38939 = net_38939;
  assign seg_10_13_neigh_op_rgt_3_42766 = seg_11_13_lutff_3_out_42766;
  assign seg_10_13_neigh_op_rgt_7_42770 = seg_11_13_lutff_7_out_42770;
  assign seg_10_13_neigh_op_top_0_39055 = seg_10_14_lutff_0_out_39055;
  assign seg_10_13_neigh_op_top_1_39056 = seg_10_14_lutff_1_out_39056;
  assign seg_10_13_neigh_op_top_3_39058 = seg_10_14_lutff_3_out_39058;
  assign seg_10_13_sp4_h_r_0_42898 = net_42898;
  assign seg_10_13_sp4_h_r_6_42906 = net_42906;
  assign seg_10_13_sp4_r_v_b_30_42794 = seg_11_15_sp4_v_b_6_42794;
  assign seg_10_13_sp4_v_b_24_38957 = seg_10_15_sp4_v_b_0_38957;
  assign seg_10_13_sp4_v_t_41_39207 = seg_10_17_sp4_v_b_4_39207;
  assign seg_10_13_sp4_v_t_43_39209 = seg_10_17_sp4_v_b_6_39209;
  assign seg_10_13_sp4_v_t_45_39211 = seg_10_17_sp4_v_b_8_39211;
  assign seg_10_13_sp4_v_t_47_39213 = seg_10_17_sp4_v_b_10_39213;
  assign seg_10_14_lutff_0_out_39055 = net_39055;
  assign seg_10_14_lutff_1_out_39056 = net_39056;
  assign seg_10_14_lutff_2_out_39057 = net_39057;
  assign seg_10_14_lutff_3_out_39058 = net_39058;
  assign seg_10_14_lutff_4_out_39059 = net_39059;
  assign seg_10_14_lutff_6_out_39061 = net_39061;
  assign seg_10_14_lutff_7_out_39062 = net_39062;
  assign seg_10_14_sp4_h_r_4_43027 = net_43027;
  assign seg_10_14_sp4_r_v_b_11_42674 = net_42674;
  assign seg_10_14_sp4_v_b_11_38843 = seg_9_12_sp4_r_v_b_35_38843;
  assign seg_10_14_sp4_v_t_36_39325 = seg_10_17_sp4_v_b_12_39325;
  assign seg_10_14_sp4_v_t_37_39326 = seg_10_18_sp4_v_b_0_39326;
  assign seg_10_14_sp4_v_t_38_39327 = seg_10_17_sp4_v_b_14_39327;
  assign seg_10_14_sp4_v_t_39_39328 = seg_10_18_sp4_v_b_2_39328;
  assign seg_10_14_sp4_v_t_41_39330 = seg_10_18_sp4_v_b_4_39330;
  assign seg_10_14_sp4_v_t_43_39332 = seg_10_18_sp4_v_b_6_39332;
  assign seg_10_14_sp4_v_t_45_39334 = seg_10_18_sp4_v_b_8_39334;
  assign seg_10_14_sp4_v_t_47_39336 = seg_10_18_sp4_v_b_10_39336;
  assign seg_10_15_lutff_2_out_39180 = net_39180;
  assign seg_10_15_sp4_h_r_4_43150 = net_43150;
  assign seg_10_15_sp4_h_r_6_43152 = seg_12_15_sp4_h_r_30_43152;
  assign seg_10_15_sp4_v_b_0_38957 = net_38957;
  assign seg_10_15_sp4_v_b_32_39211 = seg_10_17_sp4_v_b_8_39211;
  assign seg_10_15_sp4_v_b_8_38965 = net_38965;
  assign seg_10_15_sp4_v_t_36_39448 = seg_10_18_sp4_v_b_12_39448;
  assign seg_10_15_sp4_v_t_43_39455 = seg_10_17_sp4_v_b_30_39455;
  assign seg_10_16_sp4_v_t_42_39577 = seg_10_17_sp4_v_b_42_39577;
  assign seg_10_16_sp4_v_t_44_39579 = seg_10_17_sp4_v_b_44_39579;
  assign seg_10_17_lutff_2_out_39426 = net_39426;
  assign seg_10_17_lutff_3_out_39427 = net_39427;
  assign seg_10_17_lutff_4_out_39428 = net_39428;
  assign seg_10_17_lutff_5_out_39429 = net_39429;
  assign seg_10_17_lutff_6_out_39430 = net_39430;
  assign seg_10_17_lutff_7_out_39431 = net_39431;
  assign seg_10_17_neigh_op_bnr_5_43137 = seg_11_16_lutff_5_out_43137;
  assign seg_10_17_neigh_op_rgt_1_43256 = seg_11_17_lutff_1_out_43256;
  assign seg_10_17_sp4_h_l_39_28343 = seg_8_17_sp4_h_r_26_28343;
  assign seg_10_17_sp4_h_r_14_39564 = net_39564;
  assign seg_10_17_sp4_h_r_20_39570 = net_39570;
  assign seg_10_17_sp4_h_r_26_35732 = net_35732;
  assign seg_10_17_sp4_h_r_28_35734 = net_35734;
  assign seg_10_17_sp4_h_r_6_43398 = net_43398;
  assign seg_10_17_sp4_h_r_8_43400 = net_43400;
  assign seg_10_17_sp4_r_v_b_11_43043 = net_43043;
  assign seg_10_17_sp4_r_v_b_13_43157 = net_43157;
  assign seg_10_17_sp4_r_v_b_15_43159 = net_43159;
  assign seg_10_17_sp4_r_v_b_25_43279 = net_43279;
  assign seg_10_17_sp4_r_v_b_27_43281 = net_43281;
  assign seg_10_17_sp4_r_v_b_29_43283 = net_43283;
  assign seg_10_17_sp4_r_v_b_31_43285 = net_43285;
  assign seg_10_17_sp4_r_v_b_37_43403 = net_43403;
  assign seg_10_17_sp4_r_v_b_39_43405 = net_43405;
  assign seg_10_17_sp4_r_v_b_41_43407 = net_43407;
  assign seg_10_17_sp4_r_v_b_5_43037 = net_43037;
  assign seg_10_17_sp4_r_v_b_9_43041 = net_43041;
  assign seg_10_17_sp4_v_b_10_39213 = net_39213;
  assign seg_10_17_sp4_v_b_12_39325 = net_39325;
  assign seg_10_17_sp4_v_b_14_39327 = net_39327;
  assign seg_10_17_sp4_v_b_30_39455 = net_39455;
  assign seg_10_17_sp4_v_b_42_39577 = net_39577;
  assign seg_10_17_sp4_v_b_44_39579 = net_39579;
  assign seg_10_17_sp4_v_b_4_39207 = net_39207;
  assign seg_10_17_sp4_v_b_6_39209 = net_39209;
  assign seg_10_17_sp4_v_b_8_39211 = net_39211;
  assign seg_10_18_lutff_0_out_39547 = net_39547;
  assign seg_10_18_lutff_1_out_39548 = net_39548;
  assign seg_10_18_lutff_2_out_39549 = net_39549;
  assign seg_10_18_lutff_3_out_39550 = net_39550;
  assign seg_10_18_lutff_4_out_39551 = net_39551;
  assign seg_10_18_lutff_5_out_39552 = net_39552;
  assign seg_10_18_lutff_6_out_39553 = net_39553;
  assign seg_10_18_lutff_7_out_39554 = net_39554;
  assign seg_10_18_sp4_h_r_14_39687 = net_39687;
  assign seg_10_18_sp4_h_r_16_39689 = net_39689;
  assign seg_10_18_sp4_h_r_18_39691 = net_39691;
  assign seg_10_18_sp4_h_r_22_39685 = net_39685;
  assign seg_10_18_sp4_h_r_24_35851 = net_35851;
  assign seg_10_18_sp4_h_r_26_35855 = net_35855;
  assign seg_10_18_sp4_h_r_32_35861 = net_35861;
  assign seg_10_18_sp4_h_r_34_35853 = net_35853;
  assign seg_10_18_sp4_h_r_4_43519 = net_43519;
  assign seg_10_18_sp4_h_r_8_43523 = net_43523;
  assign seg_10_18_sp4_r_v_b_11_43166 = net_43166;
  assign seg_10_18_sp4_r_v_b_13_43280 = net_43280;
  assign seg_10_18_sp4_r_v_b_15_43282 = net_43282;
  assign seg_10_18_sp4_r_v_b_19_43286 = net_43286;
  assign seg_10_18_sp4_r_v_b_1_43156 = net_43156;
  assign seg_10_18_sp4_r_v_b_23_43290 = net_43290;
  assign seg_10_18_sp4_r_v_b_31_43408 = net_43408;
  assign seg_10_18_sp4_r_v_b_37_43526 = net_43526;
  assign seg_10_18_sp4_r_v_b_39_43528 = net_43528;
  assign seg_10_18_sp4_r_v_b_3_43158 = net_43158;
  assign seg_10_18_sp4_r_v_b_43_43532 = net_43532;
  assign seg_10_18_sp4_r_v_b_45_43534 = net_43534;
  assign seg_10_18_sp4_r_v_b_5_43160 = net_43160;
  assign seg_10_18_sp4_r_v_b_9_43164 = net_43164;
  assign seg_10_18_sp4_v_b_0_39326 = net_39326;
  assign seg_10_18_sp4_v_b_10_39336 = net_39336;
  assign seg_10_18_sp4_v_b_11_39335 = seg_9_18_sp4_r_v_b_11_39335;
  assign seg_10_18_sp4_v_b_12_39448 = net_39448;
  assign seg_10_18_sp4_v_b_2_39328 = net_39328;
  assign seg_10_18_sp4_v_b_4_39330 = net_39330;
  assign seg_10_18_sp4_v_b_6_39332 = net_39332;
  assign seg_10_18_sp4_v_b_8_39334 = net_39334;
  assign seg_10_19_lutff_0_out_39670 = net_39670;
  assign seg_10_19_lutff_1_out_39671 = net_39671;
  assign seg_10_19_lutff_2_out_39672 = net_39672;
  assign seg_10_19_lutff_3_out_39673 = net_39673;
  assign seg_10_19_lutff_4_out_39674 = net_39674;
  assign seg_10_19_lutff_5_out_39675 = net_39675;
  assign seg_10_19_lutff_6_out_39676 = net_39676;
  assign seg_10_19_lutff_7_out_39677 = net_39677;
  assign seg_10_19_sp4_h_r_0_43636 = net_43636;
  assign seg_10_19_sp4_h_r_10_43638 = net_43638;
  assign seg_10_19_sp4_h_r_12_39806 = net_39806;
  assign seg_10_19_sp4_h_r_14_39810 = net_39810;
  assign seg_10_19_sp4_h_r_16_39812 = net_39812;
  assign seg_10_19_sp4_h_r_20_39816 = net_39816;
  assign seg_10_19_sp4_h_r_24_35974 = net_35974;
  assign seg_10_19_sp4_h_r_28_35980 = net_35980;
  assign seg_10_19_sp4_h_r_2_43640 = net_43640;
  assign seg_10_19_sp4_h_r_34_35976 = net_35976;
  assign seg_10_19_sp4_h_r_4_43642 = net_43642;
  assign seg_10_19_sp4_h_r_6_43644 = net_43644;
  assign seg_10_19_sp4_h_r_8_43646 = net_43646;
  assign seg_10_19_sp4_r_v_b_21_43411 = net_43411;
  assign seg_10_19_sp4_r_v_b_23_43413 = net_43413;
  assign seg_10_20_lutff_0_out_39793 = net_39793;
  assign seg_10_20_lutff_1_out_39794 = net_39794;
  assign seg_10_20_lutff_2_out_39795 = net_39795;
  assign seg_10_20_lutff_3_out_39796 = net_39796;
  assign seg_10_20_sp12_h_r_12_21400 = net_21400;
  assign seg_10_20_sp4_h_r_0_43759 = net_43759;
  assign seg_10_20_sp4_h_r_22_39931 = net_39931;
  assign seg_10_20_sp4_h_r_2_43763 = net_43763;
  assign seg_10_20_sp4_h_r_4_43765 = net_43765;
  assign seg_10_20_sp4_h_r_6_43767 = net_43767;
  assign seg_10_26_lutff_7_out_40538 = net_40538;
  assign seg_10_26_sp12_v_b_20_44250 = net_44250;
  assign seg_10_27_lutff_2_out_40656 = net_40656;
  assign seg_10_27_lutff_3_out_40657 = net_40657;
  assign seg_10_27_lutff_4_out_40658 = net_40658;
  assign seg_10_27_lutff_5_out_40659 = net_40659;
  assign seg_10_27_lutff_6_out_40660 = net_40660;
  assign seg_10_27_lutff_7_out_40661 = net_40661;
  assign seg_10_27_neigh_op_lft_5_36828 = seg_9_27_lutff_5_out_36828;
  assign seg_10_27_neigh_op_lft_7_36830 = seg_9_27_lutff_7_out_36830;
  assign seg_10_27_neigh_op_top_3_40780 = seg_10_28_lutff_3_out_40780;
  assign seg_10_27_neigh_op_top_7_40784 = seg_10_28_lutff_7_out_40784;
  assign seg_10_27_sp4_v_b_36_40801 = seg_10_29_sp4_v_b_12_40801;
  assign seg_10_28_lutff_2_out_40779 = net_40779;
  assign seg_10_28_lutff_3_out_40780 = net_40780;
  assign seg_10_28_lutff_7_out_40784 = net_40784;
  assign seg_10_28_neigh_op_bnl_5_36828 = seg_9_27_lutff_5_out_36828;
  assign seg_10_28_neigh_op_bnl_7_36830 = seg_9_27_lutff_7_out_36830;
  assign seg_10_28_neigh_op_bot_4_40658 = seg_10_27_lutff_4_out_40658;
  assign seg_10_28_neigh_op_bot_6_40660 = seg_10_27_lutff_6_out_40660;
  assign seg_10_28_neigh_op_bot_7_40661 = seg_10_27_lutff_7_out_40661;
  assign seg_10_28_neigh_op_tnl_3_37072 = seg_9_29_lutff_3_out_37072;
  assign seg_10_28_neigh_op_top_6_40906 = seg_10_29_lutff_6_out_40906;
  assign seg_10_28_sp4_v_b_26_40804 = net_40804;
  assign seg_10_29_lutff_0_out_40900 = net_40900;
  assign seg_10_29_lutff_2_out_40902 = net_40902;
  assign seg_10_29_lutff_3_out_40903 = net_40903;
  assign seg_10_29_lutff_5_out_40905 = net_40905;
  assign seg_10_29_lutff_6_out_40906 = net_40906;
  assign seg_10_29_lutff_7_out_40907 = net_40907;
  assign seg_10_29_neigh_op_top_3_41026 = seg_10_30_lutff_3_out_41026;
  assign seg_10_29_neigh_op_top_4_41027 = seg_10_30_lutff_4_out_41027;
  assign seg_10_29_sp4_h_l_38_29568 = seg_9_29_sp4_h_r_38_29568;
  assign seg_10_29_sp4_v_b_12_40801 = net_40801;
  assign seg_10_2_lutff_2_out_37545 = net_37545;
  assign seg_10_2_lutff_3_out_37546 = net_37546;
  assign seg_10_2_lutff_4_out_37547 = net_37547;
  assign seg_10_2_lutff_5_out_37548 = net_37548;
  assign seg_10_2_lutff_6_out_37549 = net_37549;
  assign seg_10_2_lutff_7_out_37550 = net_37550;
  assign seg_10_2_neigh_op_lft_4_33716 = seg_9_2_lutff_4_out_33716;
  assign seg_10_2_neigh_op_top_2_37704 = seg_10_3_lutff_2_out_37704;
  assign seg_10_2_neigh_op_top_3_37705 = seg_10_3_lutff_3_out_37705;
  assign seg_10_2_neigh_op_top_4_37706 = seg_10_3_lutff_4_out_37706;
  assign seg_10_2_neigh_op_top_6_37708 = seg_10_3_lutff_6_out_37708;
  assign seg_10_30_lutff_0_out_41023 = net_41023;
  assign seg_10_30_lutff_2_out_41025 = net_41025;
  assign seg_10_30_lutff_3_out_41026 = net_41026;
  assign seg_10_30_lutff_4_out_41027 = net_41027;
  assign seg_10_30_lutff_6_out_41029 = net_41029;
  assign seg_10_30_lutff_7_out_41030 = net_41030;
  assign seg_10_30_neigh_op_bot_0_40900 = seg_10_29_lutff_0_out_40900;
  assign seg_10_30_neigh_op_bot_2_40902 = seg_10_29_lutff_2_out_40902;
  assign seg_10_30_neigh_op_bot_5_40905 = seg_10_29_lutff_5_out_40905;
  assign seg_10_30_neigh_op_lft_5_37197 = seg_9_30_lutff_5_out_37197;
  assign seg_10_30_sp12_v_b_12_44250 = seg_10_26_sp12_v_b_20_44250;
  assign seg_10_30_sp4_v_b_2_40804 = seg_10_28_sp4_v_b_26_40804;
  assign seg_10_3_lutff_2_out_37704 = net_37704;
  assign seg_10_3_lutff_3_out_37705 = net_37705;
  assign seg_10_3_lutff_4_out_37706 = net_37706;
  assign seg_10_3_lutff_6_out_37708 = net_37708;
  assign seg_10_3_lutff_7_out_37709 = net_37709;
  assign seg_10_3_neigh_op_bnl_4_33716 = seg_9_2_lutff_4_out_33716;
  assign seg_10_3_neigh_op_bot_3_37546 = seg_10_2_lutff_3_out_37546;
  assign seg_10_3_neigh_op_bot_5_37548 = seg_10_2_lutff_5_out_37548;
  assign seg_10_3_sp4_h_l_43_26919 = seg_8_3_sp4_h_r_30_26919;
  assign seg_10_4_sp4_h_l_47_27015 = seg_8_4_sp4_h_r_34_27015;
  assign seg_10_6_sp4_v_b_10_37860 = seg_9_5_sp4_r_v_b_23_37860;
  assign seg_10_7_sp4_h_r_10_42162 = net_42162;
  assign seg_10_7_sp4_r_v_b_11_41813 = net_41813;
  assign seg_10_7_sp4_r_v_b_27_42051 = net_42051;
  assign seg_10_7_sp4_v_b_10_37983 = net_37983;
  assign seg_10_8_lutff_0_out_38317 = net_38317;
  assign seg_10_8_lutff_2_out_38319 = net_38319;
  assign seg_10_8_lutff_3_out_38320 = net_38320;
  assign seg_10_8_lutff_4_out_38321 = net_38321;
  assign seg_10_8_lutff_6_out_38323 = net_38323;
  assign seg_10_8_lutff_7_out_38324 = net_38324;
  assign seg_10_8_neigh_op_bnr_0_42025 = seg_11_7_lutff_0_out_42025;
  assign seg_10_8_neigh_op_lft_5_34491 = seg_9_8_lutff_5_out_34491;
  assign seg_10_8_neigh_op_lft_6_34492 = seg_9_8_lutff_6_out_34492;
  assign seg_10_8_neigh_op_lft_7_34493 = seg_9_8_lutff_7_out_34493;
  assign seg_10_8_neigh_op_rgt_5_42153 = seg_11_8_lutff_5_out_42153;
  assign seg_10_8_neigh_op_rgt_6_42154 = seg_11_8_lutff_6_out_42154;
  assign seg_10_8_neigh_op_rgt_7_42155 = seg_11_8_lutff_7_out_42155;
  assign seg_10_8_sp4_r_v_b_35_42182 = net_42182;
  assign seg_10_8_sp4_r_v_b_36_42295 = seg_11_10_sp4_v_b_12_42295;
  assign seg_10_8_sp4_v_t_38_38589 = seg_9_12_sp4_r_v_b_3_38589;
  assign seg_10_9_sp4_h_r_11_42409 = seg_11_9_sp4_h_r_22_42409;
  assign seg_10_9_sp4_h_r_5_42413 = seg_11_9_sp4_h_r_16_42413;
  assign seg_10_9_sp4_v_b_10_38229 = seg_9_8_sp4_r_v_b_23_38229;
  assign seg_10_9_sp4_v_b_8_38227 = seg_9_8_sp4_r_v_b_21_38227;
  assign seg_11_10_lutff_4_out_42398 = net_42398;
  assign seg_11_10_lutff_5_out_42399 = net_42399;
  assign seg_11_10_lutff_6_out_42400 = net_42400;
  assign seg_11_10_lutff_7_out_42401 = net_42401;
  assign seg_11_10_neigh_op_bot_7_42278 = seg_11_9_lutff_7_out_42278;
  assign seg_11_10_sp4_h_l_36_31037 = seg_10_10_sp4_h_r_36_31037;
  assign seg_11_10_sp4_h_r_11_46363 = seg_14_10_sp4_h_r_46_46363;
  assign seg_11_10_sp4_h_r_12_42530 = net_42530;
  assign seg_11_10_sp4_h_r_14_42534 = net_42534;
  assign seg_11_10_sp4_h_r_24_38698 = net_38698;
  assign seg_11_10_sp4_h_r_26_38702 = seg_9_10_sp4_h_r_2_38702;
  assign seg_11_10_sp4_h_r_36_34868 = seg_9_10_sp4_h_r_12_34868;
  assign seg_11_10_sp4_h_r_8_46370 = net_46370;
  assign seg_11_10_sp4_r_v_b_13_46127 = net_46127;
  assign seg_11_10_sp4_r_v_b_25_46249 = net_46249;
  assign seg_11_10_sp4_r_v_b_29_46253 = net_46253;
  assign seg_11_10_sp4_r_v_b_31_46255 = net_46255;
  assign seg_11_10_sp4_r_v_b_33_46257 = net_46257;
  assign seg_11_10_sp4_r_v_b_39_46375 = net_46375;
  assign seg_11_10_sp4_r_v_b_41_46377 = net_46377;
  assign seg_11_10_sp4_r_v_b_47_46383 = net_46383;
  assign seg_11_10_sp4_r_v_b_9_46011 = net_46011;
  assign seg_11_10_sp4_v_b_11_42182 = seg_10_8_sp4_r_v_b_35_42182;
  assign seg_11_10_sp4_v_b_12_42295 = net_42295;
  assign seg_11_10_sp4_v_b_24_42419 = net_42419;
  assign seg_11_10_sp4_v_b_40_42545 = net_42545;
  assign seg_11_10_sp4_v_b_44_42549 = net_42549;
  assign seg_11_11_lutff_2_out_42519 = net_42519;
  assign seg_11_11_lutff_7_out_42524 = net_42524;
  assign seg_11_12_lutff_2_out_42642 = net_42642;
  assign seg_11_12_lutff_6_out_42646 = net_42646;
  assign seg_11_12_lutff_7_out_42647 = net_42647;
  assign seg_11_12_neigh_op_lft_1_38810 = seg_10_12_lutff_1_out_38810;
  assign seg_11_12_neigh_op_lft_5_38814 = seg_10_12_lutff_5_out_38814;
  assign seg_11_12_neigh_op_lft_7_38816 = seg_10_12_lutff_7_out_38816;
  assign seg_11_12_neigh_op_rgt_1_46472 = seg_12_12_lutff_1_out_46472;
  assign seg_11_12_neigh_op_rgt_5_46476 = seg_12_12_lutff_5_out_46476;
  assign seg_11_12_neigh_op_rgt_7_46478 = seg_12_12_lutff_7_out_46478;
  assign seg_11_12_sp4_h_r_14_42780 = net_42780;
  assign seg_11_12_sp4_h_r_20_42786 = net_42786;
  assign seg_11_12_sp4_h_r_2_46610 = net_46610;
  assign seg_11_12_sp4_h_r_6_46614 = net_46614;
  assign seg_11_12_sp4_h_r_8_46616 = net_46616;
  assign seg_11_12_sp4_r_v_b_17_46377 = seg_11_10_sp4_r_v_b_41_46377;
  assign seg_11_12_sp4_v_b_0_42419 = seg_11_10_sp4_v_b_24_42419;
  assign seg_11_13_lutff_3_out_42766 = net_42766;
  assign seg_11_13_lutff_7_out_42770 = net_42770;
  assign seg_11_13_neigh_op_bot_7_42647 = seg_11_12_lutff_7_out_42647;
  assign seg_11_13_neigh_op_lft_1_38933 = seg_10_13_lutff_1_out_38933;
  assign seg_11_13_neigh_op_lft_2_38934 = seg_10_13_lutff_2_out_38934;
  assign seg_11_13_neigh_op_lft_4_38936 = seg_10_13_lutff_4_out_38936;
  assign seg_11_13_neigh_op_lft_5_38937 = seg_10_13_lutff_5_out_38937;
  assign seg_11_13_neigh_op_lft_6_38938 = seg_10_13_lutff_6_out_38938;
  assign seg_11_13_neigh_op_lft_7_38939 = seg_10_13_lutff_7_out_38939;
  assign seg_11_13_neigh_op_rgt_1_46595 = seg_12_13_lutff_1_out_46595;
  assign seg_11_13_neigh_op_rgt_2_46596 = seg_12_13_lutff_2_out_46596;
  assign seg_11_13_neigh_op_rgt_4_46598 = seg_12_13_lutff_4_out_46598;
  assign seg_11_13_neigh_op_rgt_5_46599 = seg_12_13_lutff_5_out_46599;
  assign seg_11_13_neigh_op_rgt_6_46600 = seg_12_13_lutff_6_out_46600;
  assign seg_11_13_neigh_op_rgt_7_46601 = seg_12_13_lutff_7_out_46601;
  assign seg_11_13_sp12_h_r_2_42895 = net_42895;
  assign seg_11_13_sp4_h_r_12_42899 = net_42899;
  assign seg_11_13_sp4_h_r_20_42909 = seg_13_13_sp4_h_r_44_42909;
  assign seg_11_13_sp4_h_r_24_39067 = net_39067;
  assign seg_11_13_sp4_h_r_2_46733 = net_46733;
  assign seg_11_13_sp4_h_r_32_39077 = net_39077;
  assign seg_11_13_sp4_h_r_4_46735 = net_46735;
  assign seg_11_13_sp4_v_b_5_42545 = seg_11_10_sp4_v_b_40_42545;
  assign seg_11_13_sp4_v_b_9_42549 = seg_11_10_sp4_v_b_44_42549;
  assign seg_11_13_sp4_v_t_40_43037 = seg_10_17_sp4_r_v_b_5_43037;
  assign seg_11_13_sp4_v_t_44_43041 = seg_10_17_sp4_r_v_b_9_43041;
  assign seg_11_13_sp4_v_t_46_43043 = seg_10_17_sp4_r_v_b_11_43043;
  assign seg_11_14_lutff_0_out_42886 = net_42886;
  assign seg_11_14_lutff_2_out_42888 = net_42888;
  assign seg_11_14_lutff_3_out_42889 = net_42889;
  assign seg_11_14_lutff_4_out_42890 = net_42890;
  assign seg_11_14_lutff_6_out_42892 = net_42892;
  assign seg_11_14_neigh_op_lft_4_39059 = seg_10_14_lutff_4_out_39059;
  assign seg_11_14_neigh_op_lft_6_39061 = seg_10_14_lutff_6_out_39061;
  assign seg_11_14_neigh_op_lft_7_39062 = seg_10_14_lutff_7_out_39062;
  assign seg_11_14_sp4_h_r_14_43026 = net_43026;
  assign seg_11_14_sp4_h_r_2_46856 = net_46856;
  assign seg_11_14_sp4_r_v_b_27_46743 = net_46743;
  assign seg_11_14_sp4_v_b_0_42665 = seg_10_11_sp4_r_v_b_37_42665;
  assign seg_11_14_sp4_v_t_36_43156 = seg_10_18_sp4_r_v_b_1_43156;
  assign seg_11_14_sp4_v_t_37_43157 = seg_10_17_sp4_r_v_b_13_43157;
  assign seg_11_14_sp4_v_t_38_43158 = seg_10_18_sp4_r_v_b_3_43158;
  assign seg_11_14_sp4_v_t_39_43159 = seg_10_17_sp4_r_v_b_15_43159;
  assign seg_11_14_sp4_v_t_40_43160 = seg_10_18_sp4_r_v_b_5_43160;
  assign seg_11_14_sp4_v_t_42_43162 = seg_11_17_sp4_v_b_18_43162;
  assign seg_11_14_sp4_v_t_44_43164 = seg_10_18_sp4_r_v_b_9_43164;
  assign seg_11_14_sp4_v_t_46_43166 = seg_10_18_sp4_r_v_b_11_43166;
  assign seg_11_15_lutff_2_out_43011 = net_43011;
  assign seg_11_15_lutff_4_out_43013 = net_43013;
  assign seg_11_15_lutff_6_out_43015 = net_43015;
  assign seg_11_15_neigh_op_rgt_0_46840 = seg_12_15_lutff_0_out_46840;
  assign seg_11_15_sp4_v_b_33_43041 = seg_10_17_sp4_r_v_b_9_43041;
  assign seg_11_15_sp4_v_b_6_42794 = net_42794;
  assign seg_11_15_sp4_v_t_36_43279 = seg_10_17_sp4_r_v_b_25_43279;
  assign seg_11_15_sp4_v_t_37_43280 = seg_10_18_sp4_r_v_b_13_43280;
  assign seg_11_15_sp4_v_t_38_43281 = seg_10_17_sp4_r_v_b_27_43281;
  assign seg_11_15_sp4_v_t_40_43283 = seg_10_17_sp4_r_v_b_29_43283;
  assign seg_11_15_sp4_v_t_42_43285 = seg_10_17_sp4_r_v_b_31_43285;
  assign seg_11_15_sp4_v_t_43_43286 = seg_10_18_sp4_r_v_b_19_43286;
  assign seg_11_15_sp4_v_t_47_43290 = seg_10_18_sp4_r_v_b_23_43290;
  assign seg_11_16_lutff_5_out_43137 = net_43137;
  assign seg_11_16_sp4_h_r_10_47100 = net_47100;
  assign seg_11_16_sp4_r_v_b_11_46751 = net_46751;
  assign seg_11_16_sp4_r_v_b_43_47117 = net_47117;
  assign seg_11_16_sp4_v_t_37_43403 = seg_10_17_sp4_r_v_b_37_43403;
  assign seg_11_16_sp4_v_t_39_43405 = seg_10_17_sp4_r_v_b_39_43405;
  assign seg_11_16_sp4_v_t_41_43407 = seg_10_17_sp4_r_v_b_41_43407;
  assign seg_11_17_lutff_1_out_43256 = net_43256;
  assign seg_11_17_sp4_h_r_18_43399 = net_43399;
  assign seg_11_17_sp4_h_r_2_47225 = net_47225;
  assign seg_11_17_sp4_r_v_b_35_47120 = net_47120;
  assign seg_11_17_sp4_v_b_18_43162 = net_43162;
  assign seg_11_17_sp4_v_t_37_43526 = seg_10_18_sp4_r_v_b_37_43526;
  assign seg_11_17_sp4_v_t_39_43528 = seg_10_18_sp4_r_v_b_39_43528;
  assign seg_11_17_sp4_v_t_43_43532 = seg_10_18_sp4_r_v_b_43_43532;
  assign seg_11_17_sp4_v_t_45_43534 = seg_10_18_sp4_r_v_b_45_43534;
  assign seg_11_18_lutff_3_out_43381 = net_43381;
  assign seg_11_18_lutff_4_out_43382 = net_43382;
  assign seg_11_18_lutff_5_out_43383 = net_43383;
  assign seg_11_18_neigh_op_tnl_0_39670 = seg_10_19_lutff_0_out_39670;
  assign seg_11_18_neigh_op_tnl_5_39675 = seg_10_19_lutff_5_out_39675;
  assign seg_11_18_neigh_op_tnl_6_39676 = seg_10_19_lutff_6_out_39676;
  assign seg_11_18_sp4_h_r_26_39686 = seg_9_18_sp4_h_r_2_39686;
  assign seg_11_18_sp4_h_r_2_47348 = net_47348;
  assign seg_11_18_sp4_h_r_4_47350 = net_47350;
  assign seg_11_18_sp4_r_v_b_41_47361 = seg_12_21_sp4_v_b_4_47361;
  assign seg_11_19_lutff_2_out_43503 = net_43503;
  assign seg_11_19_lutff_6_out_43507 = net_43507;
  assign seg_11_19_neigh_op_lft_1_39671 = seg_10_19_lutff_1_out_39671;
  assign seg_11_19_neigh_op_lft_4_39674 = seg_10_19_lutff_4_out_39674;
  assign seg_11_19_neigh_op_top_1_43625 = seg_11_20_lutff_1_out_43625;
  assign seg_11_19_sp4_h_r_6_47475 = net_47475;
  assign seg_11_19_sp4_r_v_b_28_47361 = seg_12_21_sp4_v_b_4_47361;
  assign seg_11_19_sp4_v_b_2_43282 = seg_10_18_sp4_r_v_b_15_43282;
  assign seg_11_20_lutff_1_out_43625 = net_43625;
  assign seg_11_20_neigh_op_bnl_4_39674 = seg_10_19_lutff_4_out_39674;
  assign seg_11_20_neigh_op_lft_1_39794 = seg_10_20_lutff_1_out_39794;
  assign seg_11_20_neigh_op_lft_2_39795 = seg_10_20_lutff_2_out_39795;
  assign seg_11_20_sp4_h_r_12_43760 = net_43760;
  assign seg_11_20_sp4_h_r_4_47596 = net_47596;
  assign seg_11_20_sp4_v_b_10_43413 = seg_10_19_sp4_r_v_b_23_43413;
  assign seg_11_20_sp4_v_b_7_43408 = seg_10_18_sp4_r_v_b_31_43408;
  assign seg_11_20_sp4_v_b_8_43411 = seg_10_19_sp4_r_v_b_21_43411;
  assign seg_11_21_sp4_h_r_5_47720 = seg_12_21_sp4_h_r_16_47720;
  assign seg_11_22_sp4_v_t_44_44148 = seg_11_23_sp4_v_b_44_44148;
  assign seg_11_23_sp4_r_v_b_13_47726 = net_47726;
  assign seg_11_23_sp4_v_b_44_44148 = net_44148;
  assign seg_11_25_sp4_v_t_47_44520 = seg_11_29_sp4_v_b_10_44520;
  assign seg_11_29_neigh_op_lft_3_40903 = seg_10_29_lutff_3_out_40903;
  assign seg_11_29_neigh_op_lft_5_40905 = seg_10_29_lutff_5_out_40905;
  assign seg_11_29_sp4_v_b_10_44520 = net_44520;
  assign seg_11_30_neigh_op_bnl_0_40900 = seg_10_29_lutff_0_out_40900;
  assign seg_11_30_neigh_op_bnl_5_40905 = seg_10_29_lutff_5_out_40905;
  assign seg_11_30_neigh_op_lft_3_41026 = seg_10_30_lutff_3_out_41026;
  assign seg_11_30_neigh_op_lft_4_41027 = seg_10_30_lutff_4_out_41027;
  assign seg_11_30_sp4_h_r_6_48824 = net_48824;
  assign seg_11_31_span4_horz_l_14_33556 = seg_8_31_span4_horz_r_6_33556;
  assign seg_11_4_sp4_h_l_42_30307 = seg_8_4_sp4_h_r_18_30307;
  assign seg_11_7_lutff_0_out_42025 = net_42025;
  assign seg_11_7_lutff_2_out_42027 = net_42027;
  assign seg_11_7_lutff_7_out_42032 = net_42032;
  assign seg_11_7_sp4_r_v_b_17_45762 = net_45762;
  assign seg_11_7_sp4_v_b_11_41813 = seg_10_7_sp4_r_v_b_11_41813;
  assign seg_11_7_sp4_v_t_36_42295 = seg_11_10_sp4_v_b_12_42295;
  assign seg_11_8_lutff_2_out_42150 = net_42150;
  assign seg_11_8_lutff_3_out_42151 = net_42151;
  assign seg_11_8_lutff_4_out_42152 = net_42152;
  assign seg_11_8_lutff_5_out_42153 = net_42153;
  assign seg_11_8_lutff_6_out_42154 = net_42154;
  assign seg_11_8_lutff_7_out_42155 = net_42155;
  assign seg_11_8_neigh_op_bot_0_42025 = seg_11_7_lutff_0_out_42025;
  assign seg_11_8_neigh_op_lft_2_38319 = seg_10_8_lutff_2_out_38319;
  assign seg_11_8_neigh_op_lft_4_38321 = seg_10_8_lutff_4_out_38321;
  assign seg_11_8_neigh_op_lft_6_38323 = seg_10_8_lutff_6_out_38323;
  assign seg_11_8_neigh_op_rgt_1_45980 = seg_12_8_lutff_1_out_45980;
  assign seg_11_8_neigh_op_top_0_42271 = seg_11_9_lutff_0_out_42271;
  assign seg_11_8_neigh_op_top_1_42272 = seg_11_9_lutff_1_out_42272;
  assign seg_11_8_neigh_op_top_3_42274 = seg_11_9_lutff_3_out_42274;
  assign seg_11_8_sp4_h_l_37_30790 = seg_9_8_sp4_h_r_24_30790;
  assign seg_11_9_lutff_0_out_42271 = net_42271;
  assign seg_11_9_lutff_1_out_42272 = net_42272;
  assign seg_11_9_lutff_3_out_42274 = net_42274;
  assign seg_11_9_lutff_4_out_42275 = net_42275;
  assign seg_11_9_lutff_5_out_42276 = net_42276;
  assign seg_11_9_lutff_6_out_42277 = net_42277;
  assign seg_11_9_lutff_7_out_42278 = net_42278;
  assign seg_11_9_neigh_op_bnr_5_45984 = seg_12_8_lutff_5_out_45984;
  assign seg_11_9_neigh_op_bot_2_42150 = seg_11_8_lutff_2_out_42150;
  assign seg_11_9_neigh_op_bot_3_42151 = seg_11_8_lutff_3_out_42151;
  assign seg_11_9_neigh_op_bot_4_42152 = seg_11_8_lutff_4_out_42152;
  assign seg_11_9_neigh_op_top_6_42400 = seg_11_10_lutff_6_out_42400;
  assign seg_11_9_sp4_h_r_16_42413 = net_42413;
  assign seg_11_9_sp4_h_r_22_42409 = net_42409;
  assign seg_11_9_sp4_h_r_34_38577 = net_38577;
  assign seg_11_9_sp4_v_b_3_42051 = seg_10_7_sp4_r_v_b_27_42051;
  assign seg_12_10_sp4_v_b_9_46011 = seg_11_10_sp4_r_v_b_9_46011;
  assign seg_12_11_lutff_0_out_46348 = net_46348;
  assign seg_12_11_lutff_2_out_46350 = net_46350;
  assign seg_12_11_lutff_5_out_46353 = net_46353;
  assign seg_12_11_lutff_6_out_46354 = net_46354;
  assign seg_12_11_neigh_op_bnl_4_42398 = seg_11_10_lutff_4_out_42398;
  assign seg_12_11_neigh_op_lft_2_42519 = seg_11_11_lutff_2_out_42519;
  assign seg_12_11_neigh_op_lft_7_42524 = seg_11_11_lutff_7_out_42524;
  assign seg_12_11_sp12_v_t_23_50313 = seg_12_21_sp12_v_b_4_50313;
  assign seg_12_11_sp4_h_r_2_50318 = net_50318;
  assign seg_12_11_sp4_r_v_b_23_50091 = net_50091;
  assign seg_12_12_lutff_1_out_46472 = net_46472;
  assign seg_12_12_lutff_3_out_46474 = net_46474;
  assign seg_12_12_lutff_4_out_46475 = net_46475;
  assign seg_12_12_lutff_5_out_46476 = net_46476;
  assign seg_12_12_lutff_6_out_46477 = net_46477;
  assign seg_12_12_lutff_7_out_46478 = net_46478;
  assign seg_12_12_neigh_op_bnr_1_50180 = seg_13_11_lutff_1_out_50180;
  assign seg_12_12_neigh_op_bot_2_46350 = seg_12_11_lutff_2_out_46350;
  assign seg_12_12_neigh_op_bot_5_46353 = seg_12_11_lutff_5_out_46353;
  assign seg_12_12_neigh_op_rgt_4_50306 = seg_13_12_lutff_4_out_50306;
  assign seg_12_12_sp4_h_r_16_46613 = seg_14_12_sp4_h_r_40_46613;
  assign seg_12_12_sp4_h_r_18_46615 = seg_14_12_sp4_h_r_42_46615;
  assign seg_12_12_sp4_h_r_4_50443 = net_50443;
  assign seg_12_12_sp4_v_b_1_46249 = seg_11_10_sp4_r_v_b_25_46249;
  assign seg_12_12_sp4_v_b_32_46504 = seg_12_14_sp4_v_b_8_46504;
  assign seg_12_12_sp4_v_b_43_46625 = seg_12_15_sp4_v_b_6_46625;
  assign seg_12_12_sp4_v_b_5_46253 = seg_11_10_sp4_r_v_b_29_46253;
  assign seg_12_12_sp4_v_b_7_46255 = seg_11_10_sp4_r_v_b_31_46255;
  assign seg_12_12_sp4_v_t_46_46751 = seg_11_16_sp4_r_v_b_11_46751;
  assign seg_12_13_lutff_0_out_46594 = net_46594;
  assign seg_12_13_lutff_1_out_46595 = net_46595;
  assign seg_12_13_lutff_2_out_46596 = net_46596;
  assign seg_12_13_lutff_3_out_46597 = net_46597;
  assign seg_12_13_lutff_4_out_46598 = net_46598;
  assign seg_12_13_lutff_5_out_46599 = net_46599;
  assign seg_12_13_lutff_6_out_46600 = net_46600;
  assign seg_12_13_lutff_7_out_46601 = net_46601;
  assign seg_12_13_neigh_op_tnl_2_42888 = seg_11_14_lutff_2_out_42888;
  assign seg_12_13_neigh_op_tnl_3_42889 = seg_11_14_lutff_3_out_42889;
  assign seg_12_13_neigh_op_tnr_2_50550 = seg_13_14_lutff_2_out_50550;
  assign seg_12_13_neigh_op_top_1_46718 = seg_12_14_lutff_1_out_46718;
  assign seg_12_13_neigh_op_top_3_46720 = seg_12_14_lutff_3_out_46720;
  assign seg_12_13_neigh_op_top_5_46722 = seg_12_14_lutff_5_out_46722;
  assign seg_12_13_sp4_h_r_8_50570 = seg_14_13_sp4_h_r_32_50570;
  assign seg_12_13_sp4_r_v_b_27_50451 = seg_12_15_sp4_r_v_b_3_50451;
  assign seg_12_13_sp4_v_b_10_46383 = seg_11_10_sp4_r_v_b_47_46383;
  assign seg_12_13_sp4_v_b_2_46375 = seg_11_10_sp4_r_v_b_39_46375;
  assign seg_12_13_sp4_v_b_4_46377 = seg_11_10_sp4_r_v_b_41_46377;
  assign seg_12_14_lutff_0_out_46717 = net_46717;
  assign seg_12_14_lutff_1_out_46718 = net_46718;
  assign seg_12_14_lutff_3_out_46720 = net_46720;
  assign seg_12_14_lutff_4_out_46721 = net_46721;
  assign seg_12_14_lutff_5_out_46722 = net_46722;
  assign seg_12_14_neigh_op_lft_4_42890 = seg_11_14_lutff_4_out_42890;
  assign seg_12_14_neigh_op_rgt_7_50555 = seg_13_14_lutff_7_out_50555;
  assign seg_12_14_neigh_op_tnl_4_43013 = seg_11_15_lutff_4_out_43013;
  assign seg_12_14_sp4_h_r_14_46857 = net_46857;
  assign seg_12_14_sp4_h_r_28_43027 = seg_10_14_sp4_h_r_4_43027;
  assign seg_12_14_sp4_h_r_4_50689 = net_50689;
  assign seg_12_14_sp4_v_b_8_46504 = net_46504;
  assign seg_12_15_lutff_0_out_46840 = net_46840;
  assign seg_12_15_lutff_4_out_46844 = net_46844;
  assign seg_12_15_lutff_5_out_46845 = net_46845;
  assign seg_12_15_lutff_7_out_46847 = net_46847;
  assign seg_12_15_neigh_op_lft_2_43011 = seg_11_15_lutff_2_out_43011;
  assign seg_12_15_neigh_op_lft_4_43013 = seg_11_15_lutff_4_out_43013;
  assign seg_12_15_neigh_op_lft_6_43015 = seg_11_15_lutff_6_out_43015;
  assign seg_12_15_sp4_h_r_28_43150 = seg_10_15_sp4_h_r_4_43150;
  assign seg_12_15_sp4_h_r_30_43152 = net_43152;
  assign seg_12_15_sp4_h_r_4_50812 = net_50812;
  assign seg_12_15_sp4_r_v_b_3_50451 = net_50451;
  assign seg_12_15_sp4_v_b_6_46625 = net_46625;
  assign seg_12_15_sp4_v_t_43_47117 = seg_11_16_sp4_r_v_b_43_47117;
  assign seg_12_15_sp4_v_t_46_47120 = seg_11_17_sp4_r_v_b_35_47120;
  assign seg_12_16_lutff_1_out_46964 = net_46964;
  assign seg_12_16_lutff_2_out_46965 = net_46965;
  assign seg_12_16_lutff_4_out_46967 = net_46967;
  assign seg_12_16_lutff_5_out_46968 = net_46968;
  assign seg_12_16_lutff_6_out_46969 = net_46969;
  assign seg_12_16_neigh_op_top_1_47087 = seg_12_17_lutff_1_out_47087;
  assign seg_12_16_sp4_h_r_8_50939 = net_50939;
  assign seg_12_16_sp4_v_b_3_46743 = seg_11_14_sp4_r_v_b_27_46743;
  assign seg_12_17_lutff_0_out_47086 = net_47086;
  assign seg_12_17_lutff_1_out_47087 = net_47087;
  assign seg_12_17_lutff_3_out_47089 = net_47089;
  assign seg_12_17_lutff_5_out_47091 = net_47091;
  assign seg_12_17_lutff_6_out_47092 = net_47092;
  assign seg_12_17_neigh_op_bot_4_46967 = seg_12_16_lutff_4_out_46967;
  assign seg_12_17_sp4_h_l_39_35732 = seg_10_17_sp4_h_r_26_35732;
  assign seg_12_17_sp4_h_l_41_35734 = seg_10_17_sp4_h_r_28_35734;
  assign seg_12_17_sp4_h_r_10_51054 = net_51054;
  assign seg_12_17_sp4_h_r_38_39564 = seg_10_17_sp4_h_r_14_39564;
  assign seg_12_17_sp4_v_t_37_47357 = seg_12_21_sp4_v_b_0_47357;
  assign seg_12_17_sp4_v_t_41_47361 = seg_12_21_sp4_v_b_4_47361;
  assign seg_12_17_sp4_v_t_45_47365 = seg_12_21_sp4_v_b_8_47365;
  assign seg_12_18_lutff_2_out_47211 = net_47211;
  assign seg_12_18_lutff_5_out_47214 = net_47214;
  assign seg_12_18_lutff_7_out_47216 = net_47216;
  assign seg_12_18_neigh_op_lft_4_43382 = seg_11_18_lutff_4_out_43382;
  assign seg_12_18_neigh_op_rgt_4_51044 = seg_13_18_lutff_4_out_51044;
  assign seg_12_18_neigh_op_top_7_47339 = seg_12_19_lutff_7_out_47339;
  assign seg_12_18_sp4_h_l_37_35851 = seg_10_18_sp4_h_r_24_35851;
  assign seg_12_18_sp4_h_l_39_35855 = seg_10_18_sp4_h_r_26_35855;
  assign seg_12_18_sp4_h_l_45_35861 = seg_10_18_sp4_h_r_32_35861;
  assign seg_12_18_sp4_h_l_47_35853 = seg_10_18_sp4_h_r_34_35853;
  assign seg_12_18_sp4_h_r_0_51175 = net_51175;
  assign seg_12_18_sp4_h_r_16_47351 = net_47351;
  assign seg_12_18_sp4_v_b_41_47361 = seg_12_21_sp4_v_b_4_47361;
  assign seg_12_18_sp4_v_t_40_47483 = seg_12_21_sp4_v_b_16_47483;
  assign seg_12_19_lutff_3_out_47335 = net_47335;
  assign seg_12_19_lutff_4_out_47336 = net_47336;
  assign seg_12_19_lutff_6_out_47338 = net_47338;
  assign seg_12_19_lutff_7_out_47339 = net_47339;
  assign seg_12_19_neigh_op_lft_2_43503 = seg_11_19_lutff_2_out_43503;
  assign seg_12_19_neigh_op_top_1_47456 = seg_12_20_lutff_1_out_47456;
  assign seg_12_19_sp4_h_l_37_35974 = seg_10_19_sp4_h_r_24_35974;
  assign seg_12_19_sp4_h_l_41_35980 = seg_10_19_sp4_h_r_28_35980;
  assign seg_12_19_sp4_h_l_47_35976 = seg_10_19_sp4_h_r_34_35976;
  assign seg_12_19_sp4_h_r_24_43636 = seg_10_19_sp4_h_r_0_43636;
  assign seg_12_19_sp4_h_r_32_43646 = seg_10_19_sp4_h_r_8_43646;
  assign seg_12_19_sp4_h_r_3_51303 = seg_15_19_sp4_h_r_38_51303;
  assign seg_12_19_sp4_h_r_4_51304 = net_51304;
  assign seg_12_19_sp4_r_v_b_37_51311 = net_51311;
  assign seg_12_19_sp4_v_t_37_47603 = seg_12_23_sp4_v_b_0_47603;
  assign seg_12_20_lutff_1_out_47456 = net_47456;
  assign seg_12_21_lutff_2_out_47580 = net_47580;
  assign seg_12_21_lutff_6_out_47584 = net_47584;
  assign seg_12_21_neigh_op_tnr_3_51535 = seg_13_22_lutff_3_out_51535;
  assign seg_12_21_neigh_op_tnr_7_51539 = seg_13_22_lutff_7_out_51539;
  assign seg_12_21_sp12_v_b_4_50313 = net_50313;
  assign seg_12_21_sp12_v_t_23_51543 = seg_12_31_span12_vert_4_51543;
  assign seg_12_21_sp4_h_r_0_51544 = net_51544;
  assign seg_12_21_sp4_h_r_14_47718 = net_47718;
  assign seg_12_21_sp4_h_r_16_47720 = net_47720;
  assign seg_12_21_sp4_h_r_20_47724 = net_47724;
  assign seg_12_21_sp4_h_r_32_43892 = net_43892;
  assign seg_12_21_sp4_h_r_4_51550 = net_51550;
  assign seg_12_21_sp4_h_r_9_51555 = seg_15_21_sp4_h_r_44_51555;
  assign seg_12_21_sp4_r_v_b_17_51315 = net_51315;
  assign seg_12_21_sp4_r_v_b_1_51187 = net_51187;
  assign seg_12_21_sp4_r_v_b_21_51319 = net_51319;
  assign seg_12_21_sp4_r_v_b_5_51191 = net_51191;
  assign seg_12_21_sp4_r_v_b_9_51195 = net_51195;
  assign seg_12_21_sp4_v_b_0_47357 = net_47357;
  assign seg_12_21_sp4_v_b_16_47483 = net_47483;
  assign seg_12_21_sp4_v_b_37_47726 = seg_11_23_sp4_r_v_b_13_47726;
  assign seg_12_21_sp4_v_b_4_47361 = net_47361;
  assign seg_12_21_sp4_v_b_8_47365 = net_47365;
  assign seg_12_23_sp4_h_r_32_44138 = net_44138;
  assign seg_12_23_sp4_r_v_b_1_51433 = net_51433;
  assign seg_12_23_sp4_v_b_0_47603 = net_47603;
  assign seg_12_27_lutff_2_out_48318 = net_48318;
  assign seg_12_27_lutff_3_out_48319 = net_48319;
  assign seg_12_27_lutff_4_out_48320 = net_48320;
  assign seg_12_27_lutff_5_out_48321 = net_48321;
  assign seg_12_27_lutff_6_out_48322 = net_48322;
  assign seg_12_27_lutff_7_out_48323 = net_48323;
  assign seg_12_27_neigh_op_rgt_4_52151 = seg_13_27_lutff_4_out_52151;
  assign seg_12_27_neigh_op_rgt_5_52152 = seg_13_27_lutff_5_out_52152;
  assign seg_12_27_neigh_op_rgt_7_52154 = seg_13_27_lutff_7_out_52154;
  assign seg_12_27_neigh_op_top_1_48440 = seg_12_28_lutff_1_out_48440;
  assign seg_12_27_sp4_h_r_12_48452 = net_48452;
  assign seg_12_27_sp4_h_r_14_48456 = net_48456;
  assign seg_12_28_lutff_1_out_48440 = net_48440;
  assign seg_12_28_lutff_2_out_48441 = net_48441;
  assign seg_12_28_sp4_h_r_10_52407 = seg_14_28_sp4_h_r_34_52407;
  assign seg_12_28_sp4_h_r_11_52408 = seg_15_28_sp4_h_r_46_52408;
  assign seg_12_28_sp4_h_r_18_48583 = net_48583;
  assign seg_12_31_span12_vert_4_51543 = net_51543;
  assign seg_12_4_sp4_h_l_39_34133 = seg_8_4_sp4_h_r_2_34133;
  assign seg_12_7_sp4_v_t_37_46127 = seg_11_10_sp4_r_v_b_13_46127;
  assign seg_12_8_lutff_1_out_45980 = net_45980;
  assign seg_12_8_lutff_5_out_45984 = net_45984;
  assign seg_12_8_neigh_op_bnl_0_42025 = seg_11_7_lutff_0_out_42025;
  assign seg_12_8_sp4_h_r_2_49949 = net_49949;
  assign seg_12_8_sp4_h_r_44_38463 = net_38463;
  assign seg_12_8_sp4_v_b_37_46127 = seg_11_10_sp4_r_v_b_13_46127;
  assign seg_12_8_sp4_v_b_4_45762 = seg_11_7_sp4_r_v_b_17_45762;
  assign seg_13_10_sp4_h_l_37_38698 = seg_11_10_sp4_h_r_24_38698;
  assign seg_13_10_sp4_h_r_0_54022 = seg_15_10_sp4_h_r_24_54022;
  assign seg_13_11_lutff_1_out_50180 = net_50180;
  assign seg_13_11_lutff_6_out_50185 = net_50185;
  assign seg_13_11_sp4_h_l_47_38823 = seg_9_11_sp4_h_r_10_38823;
  assign seg_13_12_lutff_1_out_50303 = net_50303;
  assign seg_13_12_lutff_2_out_50304 = net_50304;
  assign seg_13_12_lutff_4_out_50306 = net_50306;
  assign seg_13_12_lutff_5_out_50307 = net_50307;
  assign seg_13_12_neigh_op_lft_3_46474 = seg_12_12_lutff_3_out_46474;
  assign seg_13_12_neigh_op_lft_4_46475 = seg_12_12_lutff_4_out_46475;
  assign seg_13_12_neigh_op_lft_6_46477 = seg_12_12_lutff_6_out_46477;
  assign seg_13_12_neigh_op_top_4_50429 = seg_13_13_lutff_4_out_50429;
  assign seg_13_12_sp4_h_l_36_38945 = seg_10_12_sp4_h_r_12_38945;
  assign seg_13_12_sp4_h_r_0_54268 = net_54268;
  assign seg_13_12_sp4_h_r_28_46612 = net_46612;
  assign seg_13_12_sp4_h_r_41_42781 = seg_10_12_sp4_h_r_4_42781;
  assign seg_13_12_sp4_h_r_43_42783 = seg_10_12_sp4_h_r_6_42783;
  assign seg_13_12_sp4_h_r_44_42786 = seg_11_12_sp4_h_r_20_42786;
  assign seg_13_12_sp4_h_r_45_42785 = seg_10_12_sp4_h_r_8_42785;
  assign seg_13_12_sp4_h_r_46_42778 = net_42778;
  assign seg_13_12_sp4_h_r_5_54275 = seg_16_12_sp4_h_r_40_54275;
  assign seg_13_12_sp4_h_r_6_54276 = net_54276;
  assign seg_13_12_sp4_v_b_10_50091 = seg_12_11_sp4_r_v_b_23_50091;
  assign seg_13_13_lutff_3_out_50428 = net_50428;
  assign seg_13_13_lutff_4_out_50429 = net_50429;
  assign seg_13_13_lutff_5_out_50430 = net_50430;
  assign seg_13_13_lutff_6_out_50431 = net_50431;
  assign seg_13_13_neigh_op_bot_2_50304 = seg_13_12_lutff_2_out_50304;
  assign seg_13_13_neigh_op_lft_0_46594 = seg_12_13_lutff_0_out_46594;
  assign seg_13_13_neigh_op_lft_3_46597 = seg_12_13_lutff_3_out_46597;
  assign seg_13_13_neigh_op_top_4_50552 = seg_13_14_lutff_4_out_50552;
  assign seg_13_13_sp4_h_l_37_39067 = seg_11_13_sp4_h_r_24_39067;
  assign seg_13_13_sp4_h_l_45_39077 = seg_11_13_sp4_h_r_32_39077;
  assign seg_13_13_sp4_h_r_16_50567 = net_50567;
  assign seg_13_13_sp4_h_r_2_54395 = net_54395;
  assign seg_13_13_sp4_h_r_30_46737 = net_46737;
  assign seg_13_13_sp4_h_r_37_42898 = seg_10_13_sp4_h_r_0_42898;
  assign seg_13_13_sp4_h_r_43_42906 = seg_10_13_sp4_h_r_6_42906;
  assign seg_13_13_sp4_h_r_44_42909 = net_42909;
  assign seg_13_13_sp4_h_r_4_54397 = net_54397;
  assign seg_13_13_sp4_r_v_b_17_54162 = net_54162;
  assign seg_13_14_lutff_2_out_50550 = net_50550;
  assign seg_13_14_lutff_3_out_50551 = net_50551;
  assign seg_13_14_lutff_4_out_50552 = net_50552;
  assign seg_13_14_lutff_5_out_50553 = net_50553;
  assign seg_13_14_lutff_7_out_50555 = net_50555;
  assign seg_13_14_neigh_op_bot_5_50430 = seg_13_13_lutff_5_out_50430;
  assign seg_13_14_neigh_op_bot_6_50431 = seg_13_13_lutff_6_out_50431;
  assign seg_13_14_sp4_h_r_0_54514 = net_54514;
  assign seg_13_14_sp4_r_v_b_13_54281 = net_54281;
  assign seg_13_14_sp4_r_v_b_31_54409 = seg_13_16_sp4_r_v_b_7_54409;
  assign seg_13_14_sp4_r_v_b_3_54159 = net_54159;
  assign seg_13_14_sp4_v_b_38_50697 = seg_13_16_sp4_v_b_14_50697;
  assign seg_13_15_lutff_1_out_50672 = net_50672;
  assign seg_13_15_lutff_2_out_50673 = net_50673;
  assign seg_13_15_lutff_4_out_50675 = net_50675;
  assign seg_13_15_lutff_6_out_50677 = net_50677;
  assign seg_13_15_neigh_op_lft_4_46844 = seg_12_15_lutff_4_out_46844;
  assign seg_13_15_neigh_op_lft_5_46845 = seg_12_15_lutff_5_out_46845;
  assign seg_13_15_neigh_op_rgt_2_54504 = seg_14_15_lutff_2_out_54504;
  assign seg_13_15_neigh_op_rgt_6_54508 = seg_14_15_lutff_6_out_54508;
  assign seg_13_15_neigh_op_tnl_5_46968 = seg_12_16_lutff_5_out_46968;
  assign seg_13_15_neigh_op_tnl_6_46969 = seg_12_16_lutff_6_out_46969;
  assign seg_13_15_sp4_h_r_0_54637 = net_54637;
  assign seg_13_15_sp4_h_r_14_50811 = net_50811;
  assign seg_13_15_sp4_h_r_16_50813 = net_50813;
  assign seg_13_15_sp4_h_r_26_46979 = net_46979;
  assign seg_13_15_sp4_h_r_2_54641 = net_54641;
  assign seg_13_15_sp4_r_v_b_23_54414 = net_54414;
  assign seg_13_15_sp4_v_b_26_50698 = seg_13_17_sp4_v_b_2_50698;
  assign seg_13_16_lutff_1_out_50795 = net_50795;
  assign seg_13_16_neigh_op_bot_4_50675 = seg_13_15_lutff_4_out_50675;
  assign seg_13_16_neigh_op_bot_6_50677 = seg_13_15_lutff_6_out_50677;
  assign seg_13_16_neigh_op_rgt_0_54625 = seg_14_16_lutff_0_out_54625;
  assign seg_13_16_neigh_op_rgt_3_54628 = seg_14_16_lutff_3_out_54628;
  assign seg_13_16_neigh_op_rgt_6_54631 = seg_14_16_lutff_6_out_54631;
  assign seg_13_16_neigh_op_rgt_7_54632 = seg_14_16_lutff_7_out_54632;
  assign seg_13_16_sp4_h_r_26_47102 = net_47102;
  assign seg_13_16_sp4_h_r_2_54764 = seg_15_16_sp4_h_r_26_54764;
  assign seg_13_16_sp4_h_r_34_47100 = seg_11_16_sp4_h_r_10_47100;
  assign seg_13_16_sp4_r_v_b_13_54527 = net_54527;
  assign seg_13_16_sp4_r_v_b_41_54777 = net_54777;
  assign seg_13_16_sp4_r_v_b_5_54407 = net_54407;
  assign seg_13_16_sp4_r_v_b_7_54409 = net_54409;
  assign seg_13_16_sp4_v_b_14_50697 = net_50697;
  assign seg_13_16_sp4_v_t_43_51071 = seg_13_20_sp4_v_b_6_51071;
  assign seg_13_17_lutff_6_out_50923 = net_50923;
  assign seg_13_17_neigh_op_bnl_1_46964 = seg_12_16_lutff_1_out_46964;
  assign seg_13_17_neigh_op_lft_0_47086 = seg_12_17_lutff_0_out_47086;
  assign seg_13_17_neigh_op_lft_3_47089 = seg_12_17_lutff_3_out_47089;
  assign seg_13_17_neigh_op_lft_6_47092 = seg_12_17_lutff_6_out_47092;
  assign seg_13_17_neigh_op_rgt_2_54750 = seg_14_17_lutff_2_out_54750;
  assign seg_13_17_neigh_op_rgt_3_54751 = seg_14_17_lutff_3_out_54751;
  assign seg_13_17_neigh_op_rgt_7_54755 = seg_14_17_lutff_7_out_54755;
  assign seg_13_17_sp4_h_l_38_39564 = seg_10_17_sp4_h_r_14_39564;
  assign seg_13_17_sp4_h_l_44_39570 = seg_10_17_sp4_h_r_20_39570;
  assign seg_13_17_sp4_h_r_16_51059 = net_51059;
  assign seg_13_17_sp4_h_r_20_51063 = net_51063;
  assign seg_13_17_sp4_h_r_22_51055 = net_51055;
  assign seg_13_17_sp4_h_r_4_54889 = seg_15_17_sp4_h_r_28_54889;
  assign seg_13_17_sp4_r_v_b_11_54536 = net_54536;
  assign seg_13_17_sp4_r_v_b_15_54652 = net_54652;
  assign seg_13_17_sp4_r_v_b_41_54900 = net_54900;
  assign seg_13_17_sp4_v_b_2_50698 = net_50698;
  assign seg_13_17_sp4_v_t_36_51187 = seg_12_21_sp4_r_v_b_1_51187;
  assign seg_13_17_sp4_v_t_40_51191 = seg_12_21_sp4_r_v_b_5_51191;
  assign seg_13_17_sp4_v_t_44_51195 = seg_12_21_sp4_r_v_b_9_51195;
  assign seg_13_18_lutff_3_out_51043 = net_51043;
  assign seg_13_18_lutff_4_out_51044 = net_51044;
  assign seg_13_18_lutff_5_out_51045 = net_51045;
  assign seg_13_18_sp4_h_l_38_39687 = seg_10_18_sp4_h_r_14_39687;
  assign seg_13_18_sp4_h_l_40_39689 = seg_10_18_sp4_h_r_16_39689;
  assign seg_13_18_sp4_h_l_42_39691 = seg_10_18_sp4_h_r_18_39691;
  assign seg_13_18_sp4_h_l_46_39685 = seg_10_18_sp4_h_r_22_39685;
  assign seg_13_18_sp4_v_t_36_51310 = seg_13_21_sp4_v_b_12_51310;
  assign seg_13_18_sp4_v_t_37_51311 = seg_12_19_sp4_r_v_b_37_51311;
  assign seg_13_18_sp4_v_t_41_51315 = seg_12_21_sp4_r_v_b_17_51315;
  assign seg_13_18_sp4_v_t_45_51319 = seg_12_21_sp4_r_v_b_21_51319;
  assign seg_13_19_lutff_2_out_51165 = net_51165;
  assign seg_13_19_lutff_6_out_51169 = net_51169;
  assign seg_13_19_lutff_7_out_51170 = net_51170;
  assign seg_13_19_neigh_op_bnl_7_47216 = seg_12_18_lutff_7_out_47216;
  assign seg_13_19_neigh_op_rgt_6_55000 = seg_14_19_lutff_6_out_55000;
  assign seg_13_19_neigh_op_rgt_7_55001 = seg_14_19_lutff_7_out_55001;
  assign seg_13_19_neigh_op_top_0_51286 = seg_13_20_lutff_0_out_51286;
  assign seg_13_19_neigh_op_top_7_51293 = seg_13_20_lutff_7_out_51293;
  assign seg_13_19_sp4_h_l_36_39806 = seg_10_19_sp4_h_r_12_39806;
  assign seg_13_19_sp4_h_l_38_39810 = seg_10_19_sp4_h_r_14_39810;
  assign seg_13_19_sp4_h_l_40_39812 = seg_10_19_sp4_h_r_16_39812;
  assign seg_13_19_sp4_h_l_44_39816 = seg_10_19_sp4_h_r_20_39816;
  assign seg_13_19_sp4_h_r_18_51307 = net_51307;
  assign seg_13_19_sp4_h_r_2_55133 = net_55133;
  assign seg_13_19_sp4_h_r_41_43642 = seg_10_19_sp4_h_r_4_43642;
  assign seg_13_19_sp4_h_r_8_55139 = net_55139;
  assign seg_13_19_sp4_r_v_b_25_55018 = net_55018;
  assign seg_13_19_sp4_v_b_29_51191 = seg_12_21_sp4_r_v_b_5_51191;
  assign seg_13_19_sp4_v_t_36_51433 = seg_12_23_sp4_r_v_b_1_51433;
  assign seg_13_20_lutff_0_out_51286 = net_51286;
  assign seg_13_20_lutff_1_out_51287 = net_51287;
  assign seg_13_20_lutff_4_out_51290 = net_51290;
  assign seg_13_20_lutff_5_out_51291 = net_51291;
  assign seg_13_20_lutff_6_out_51292 = net_51292;
  assign seg_13_20_lutff_7_out_51293 = net_51293;
  assign seg_13_20_neigh_op_tnl_2_47580 = seg_12_21_lutff_2_out_47580;
  assign seg_13_20_sp12_v_b_23_55128 = seg_13_31_span12_vert_0_55128;
  assign seg_13_20_sp4_h_l_46_39931 = seg_10_20_sp4_h_r_22_39931;
  assign seg_13_20_sp4_h_r_28_47596 = seg_11_20_sp4_h_r_4_47596;
  assign seg_13_20_sp4_h_r_36_43760 = seg_11_20_sp4_h_r_12_43760;
  assign seg_13_20_sp4_h_r_37_43759 = seg_10_20_sp4_h_r_0_43759;
  assign seg_13_20_sp4_h_r_39_43763 = seg_10_20_sp4_h_r_2_43763;
  assign seg_13_20_sp4_h_r_41_43765 = seg_10_20_sp4_h_r_4_43765;
  assign seg_13_20_sp4_h_r_6_55260 = seg_15_20_sp4_h_r_30_55260;
  assign seg_13_20_sp4_v_b_6_51071 = net_51071;
  assign seg_13_21_lutff_6_out_51415 = net_51415;
  assign seg_13_21_sp12_v_b_20_55128 = seg_13_31_span12_vert_0_55128;
  assign seg_13_21_sp4_v_b_12_51310 = net_51310;
  assign seg_13_21_sp4_v_b_1_51187 = seg_12_21_sp4_r_v_b_1_51187;
  assign seg_13_21_sp4_v_t_38_51681 = seg_13_22_sp4_v_b_38_51681;
  assign seg_13_22_lutff_1_out_51533 = net_51533;
  assign seg_13_22_lutff_3_out_51535 = net_51535;
  assign seg_13_22_lutff_5_out_51537 = net_51537;
  assign seg_13_22_lutff_7_out_51539 = net_51539;
  assign seg_13_22_neigh_op_bot_6_51415 = seg_13_21_lutff_6_out_51415;
  assign seg_13_22_sp12_v_b_19_55128 = seg_13_31_span12_vert_0_55128;
  assign seg_13_22_sp12_v_b_21_55250 = seg_13_31_span12_vert_2_55250;
  assign seg_13_22_sp4_v_b_38_51681 = net_51681;
  assign seg_13_27_lutff_2_out_52149 = net_52149;
  assign seg_13_27_lutff_4_out_52151 = net_52151;
  assign seg_13_27_lutff_5_out_52152 = net_52152;
  assign seg_13_27_lutff_7_out_52154 = net_52154;
  assign seg_13_27_neigh_op_lft_4_48320 = seg_12_27_lutff_4_out_48320;
  assign seg_13_27_neigh_op_lft_5_48321 = seg_12_27_lutff_5_out_48321;
  assign seg_13_27_neigh_op_lft_6_48322 = seg_12_27_lutff_6_out_48322;
  assign seg_13_27_neigh_op_lft_7_48323 = seg_12_27_lutff_7_out_48323;
  assign seg_13_27_neigh_op_tnl_1_48440 = seg_12_28_lutff_1_out_48440;
  assign seg_13_27_sp4_r_v_b_13_55880 = net_55880;
  assign seg_13_28_sp4_h_r_6_56244 = seg_15_28_sp4_h_r_30_56244;
  assign seg_13_28_sp4_h_r_7_56245 = seg_14_28_sp4_h_r_18_56245;
  assign seg_13_31_span12_vert_0_55128 = net_55128;
  assign seg_13_31_span12_vert_2_55250 = net_55250;
  assign seg_13_3_lutff_7_out_49202 = net_49202;
  assign seg_13_3_neigh_op_tnr_1_53150 = seg_14_4_lutff_1_out_53150;
  assign seg_13_3_neigh_op_tnr_4_53153 = seg_14_4_lutff_4_out_53153;
  assign seg_13_3_neigh_op_top_6_49324 = seg_13_4_lutff_6_out_49324;
  assign seg_13_3_neigh_op_top_7_49325 = seg_13_4_lutff_7_out_49325;
  assign seg_13_3_sp4_r_v_b_19_52929 = net_52929;
  assign seg_13_4_lutff_2_out_49320 = net_49320;
  assign seg_13_4_lutff_3_out_49321 = net_49321;
  assign seg_13_4_lutff_4_out_49322 = net_49322;
  assign seg_13_4_lutff_5_out_49323 = net_49323;
  assign seg_13_4_lutff_6_out_49324 = net_49324;
  assign seg_13_4_lutff_7_out_49325 = net_49325;
  assign seg_13_4_neigh_op_bnr_0_53026 = seg_14_3_lutff_0_out_53026;
  assign seg_13_4_neigh_op_rgt_0_53149 = seg_14_4_lutff_0_out_53149;
  assign seg_13_4_neigh_op_rgt_1_53150 = seg_14_4_lutff_1_out_53150;
  assign seg_13_4_neigh_op_rgt_2_53151 = seg_14_4_lutff_2_out_53151;
  assign seg_13_4_neigh_op_rgt_4_53153 = seg_14_4_lutff_4_out_53153;
  assign seg_13_4_neigh_op_rgt_7_53156 = seg_14_4_lutff_7_out_53156;
  assign seg_13_8_lutff_2_out_49812 = net_49812;
  assign seg_13_8_lutff_3_out_49813 = net_49813;
  assign seg_13_8_lutff_4_out_49814 = net_49814;
  assign seg_13_8_lutff_5_out_49815 = net_49815;
  assign seg_13_8_lutff_7_out_49817 = net_49817;
  assign seg_13_8_neigh_op_bnr_6_53524 = seg_14_7_lutff_6_out_53524;
  assign seg_13_8_neigh_op_rgt_6_53647 = seg_14_8_lutff_6_out_53647;
  assign seg_13_8_neigh_op_rgt_7_53648 = seg_14_8_lutff_7_out_53648;
  assign seg_13_8_neigh_op_top_0_49933 = seg_13_9_lutff_0_out_49933;
  assign seg_13_8_neigh_op_top_1_49934 = seg_13_9_lutff_1_out_49934;
  assign seg_13_8_neigh_op_top_5_49938 = seg_13_9_lutff_5_out_49938;
  assign seg_13_8_neigh_op_top_6_49939 = seg_13_9_lutff_6_out_49939;
  assign seg_13_8_sp4_h_l_44_38463 = seg_12_8_sp4_h_r_44_38463;
  assign seg_13_8_sp4_h_r_12_49946 = net_49946;
  assign seg_13_8_sp4_h_r_8_53786 = seg_15_8_sp4_h_r_32_53786;
  assign seg_13_9_lutff_0_out_49933 = net_49933;
  assign seg_13_9_lutff_1_out_49934 = net_49934;
  assign seg_13_9_lutff_5_out_49938 = net_49938;
  assign seg_13_9_lutff_6_out_49939 = net_49939;
  assign seg_13_9_neigh_op_bnr_6_53647 = seg_14_8_lutff_6_out_53647;
  assign seg_13_9_neigh_op_bot_2_49812 = seg_13_8_lutff_2_out_49812;
  assign seg_13_9_neigh_op_bot_4_49814 = seg_13_8_lutff_4_out_49814;
  assign seg_13_9_neigh_op_bot_5_49815 = seg_13_8_lutff_5_out_49815;
  assign seg_13_9_neigh_op_bot_7_49817 = seg_13_8_lutff_7_out_49817;
  assign seg_13_9_neigh_op_rgt_2_53766 = seg_14_9_lutff_2_out_53766;
  assign seg_13_9_neigh_op_rgt_4_53768 = seg_14_9_lutff_4_out_53768;
  assign seg_13_9_neigh_op_rgt_5_53769 = seg_14_9_lutff_5_out_53769;
  assign seg_13_9_neigh_op_rgt_7_53771 = seg_14_9_lutff_7_out_53771;
  assign seg_13_9_sp4_r_v_b_21_53674 = net_53674;
  assign seg_14_10_neigh_op_bnr_5_57599 = seg_15_9_lutff_5_out_57599;
  assign seg_14_10_sp4_h_l_36_42530 = seg_11_10_sp4_h_r_12_42530;
  assign seg_14_10_sp4_h_l_38_42534 = seg_11_10_sp4_h_r_14_42534;
  assign seg_14_10_sp4_h_r_45_46370 = seg_11_10_sp4_h_r_8_46370;
  assign seg_14_10_sp4_h_r_46_46363 = net_46363;
  assign seg_14_10_sp4_v_b_8_53674 = seg_13_9_sp4_r_v_b_21_53674;
  assign seg_14_11_lutff_0_out_54010 = net_54010;
  assign seg_14_11_lutff_1_out_54011 = net_54011;
  assign seg_14_11_lutff_3_out_54013 = net_54013;
  assign seg_14_11_lutff_5_out_54015 = net_54015;
  assign seg_14_11_lutff_6_out_54016 = net_54016;
  assign seg_14_11_lutff_7_out_54017 = net_54017;
  assign seg_14_11_neigh_op_bnr_4_57721 = seg_15_10_lutff_4_out_57721;
  assign seg_14_11_neigh_op_lft_6_50185 = seg_13_11_lutff_6_out_50185;
  assign seg_14_11_sp4_h_r_11_57978 = seg_15_11_sp4_h_r_22_57978;
  assign seg_14_11_sp4_h_r_26_50318 = seg_12_11_sp4_h_r_2_50318;
  assign seg_14_11_sp4_h_r_4_57981 = net_57981;
  assign seg_14_11_sp4_r_v_b_37_57988 = net_57988;
  assign seg_14_11_sp4_v_b_40_54161 = net_54161;
  assign seg_14_11_sp4_v_b_45_54166 = seg_14_14_sp4_v_b_8_54166;
  assign seg_14_12_lutff_1_out_54134 = net_54134;
  assign seg_14_12_lutff_2_out_54135 = net_54135;
  assign seg_14_12_lutff_3_out_54136 = net_54136;
  assign seg_14_12_lutff_6_out_54139 = net_54139;
  assign seg_14_12_neigh_op_bnr_1_57841 = seg_15_11_lutff_1_out_57841;
  assign seg_14_12_neigh_op_bnr_2_57842 = seg_15_11_lutff_2_out_57842;
  assign seg_14_12_neigh_op_bnr_7_57847 = seg_15_11_lutff_7_out_57847;
  assign seg_14_12_neigh_op_bot_3_54013 = seg_14_11_lutff_3_out_54013;
  assign seg_14_12_sp4_h_l_38_42780 = seg_11_12_sp4_h_r_14_42780;
  assign seg_14_12_sp4_h_r_28_50443 = seg_12_12_sp4_h_r_4_50443;
  assign seg_14_12_sp4_h_r_2_58102 = net_58102;
  assign seg_14_12_sp4_h_r_39_46610 = seg_11_12_sp4_h_r_2_46610;
  assign seg_14_12_sp4_h_r_40_46613 = net_46613;
  assign seg_14_12_sp4_h_r_42_46615 = net_46615;
  assign seg_14_12_sp4_h_r_43_46614 = seg_11_12_sp4_h_r_6_46614;
  assign seg_14_12_sp4_r_v_b_0_57742 = seg_15_10_sp4_v_b_24_57742;
  assign seg_14_12_sp4_r_v_b_15_57867 = net_57867;
  assign seg_14_12_sp4_r_v_b_31_57993 = net_57993;
  assign seg_14_12_sp4_r_v_b_33_57995 = net_57995;
  assign seg_14_12_sp4_v_b_27_54159 = seg_13_14_sp4_r_v_b_3_54159;
  assign seg_14_12_sp4_v_b_39_54283 = seg_14_15_sp4_v_b_2_54283;
  assign seg_14_13_lutff_2_out_54258 = net_54258;
  assign seg_14_13_lutff_7_out_54263 = net_54263;
  assign seg_14_13_neigh_op_bnl_1_50303 = seg_13_12_lutff_1_out_50303;
  assign seg_14_13_neigh_op_bnr_1_57964 = seg_15_12_lutff_1_out_57964;
  assign seg_14_13_neigh_op_bnr_6_57969 = seg_15_12_lutff_6_out_57969;
  assign seg_14_13_neigh_op_bnr_7_57970 = seg_15_12_lutff_7_out_57970;
  assign seg_14_13_neigh_op_bot_2_54135 = seg_14_12_lutff_2_out_54135;
  assign seg_14_13_neigh_op_bot_3_54136 = seg_14_12_lutff_3_out_54136;
  assign seg_14_13_neigh_op_lft_3_50428 = seg_13_13_lutff_3_out_50428;
  assign seg_14_13_sp12_h_r_9_42895 = seg_11_13_sp12_h_r_2_42895;
  assign seg_14_13_sp4_h_l_36_42899 = seg_11_13_sp4_h_r_12_42899;
  assign seg_14_13_sp4_h_r_10_58223 = net_58223;
  assign seg_14_13_sp4_h_r_24_50560 = net_50560;
  assign seg_14_13_sp4_h_r_26_50564 = net_50564;
  assign seg_14_13_sp4_h_r_2_58225 = net_58225;
  assign seg_14_13_sp4_h_r_30_50568 = net_50568;
  assign seg_14_13_sp4_h_r_32_50570 = net_50570;
  assign seg_14_13_sp4_h_r_39_46733 = seg_11_13_sp4_h_r_2_46733;
  assign seg_14_13_sp4_h_r_41_46735 = seg_11_13_sp4_h_r_4_46735;
  assign seg_14_13_sp4_h_r_6_58229 = net_58229;
  assign seg_14_13_sp4_h_r_8_58231 = net_58231;
  assign seg_14_13_sp4_r_v_b_39_58236 = net_58236;
  assign seg_14_13_sp4_r_v_b_5_57868 = seg_15_10_sp4_v_b_40_57868;
  assign seg_14_13_sp4_v_b_12_54157 = net_54157;
  assign seg_14_13_sp4_v_b_28_54285 = seg_14_15_sp4_v_b_4_54285;
  assign seg_14_13_sp4_v_b_34_54291 = seg_14_15_sp4_v_b_10_54291;
  assign seg_14_13_sp4_v_b_40_54407 = seg_13_16_sp4_r_v_b_5_54407;
  assign seg_14_13_sp4_v_b_45_54412 = seg_14_16_sp4_v_b_8_54412;
  assign seg_14_13_sp4_v_b_47_54414 = seg_13_15_sp4_r_v_b_23_54414;
  assign seg_14_13_sp4_v_t_37_54527 = seg_13_16_sp4_r_v_b_13_54527;
  assign seg_14_14_lutff_1_out_54380 = net_54380;
  assign seg_14_14_lutff_5_out_54384 = net_54384;
  assign seg_14_14_lutff_6_out_54385 = net_54385;
  assign seg_14_14_neigh_op_lft_3_50551 = seg_13_14_lutff_3_out_50551;
  assign seg_14_14_neigh_op_top_0_54502 = seg_14_15_lutff_0_out_54502;
  assign seg_14_14_neigh_op_top_4_54506 = seg_14_15_lutff_4_out_54506;
  assign seg_14_14_sp4_h_l_38_43026 = seg_11_14_sp4_h_r_14_43026;
  assign seg_14_14_sp4_h_r_0_58344 = net_58344;
  assign seg_14_14_sp4_h_r_14_54519 = net_54519;
  assign seg_14_14_sp4_h_r_20_54525 = net_54525;
  assign seg_14_14_sp4_h_r_39_46856 = seg_11_14_sp4_h_r_2_46856;
  assign seg_14_14_sp4_r_v_b_23_58121 = net_58121;
  assign seg_14_14_sp4_r_v_b_33_58241 = net_58241;
  assign seg_14_14_sp4_v_b_14_54282 = net_54282;
  assign seg_14_14_sp4_v_b_1_54157 = seg_14_13_sp4_v_b_12_54157;
  assign seg_14_14_sp4_v_b_20_54288 = net_54288;
  assign seg_14_14_sp4_v_b_26_54406 = seg_14_16_sp4_v_b_2_54406;
  assign seg_14_14_sp4_v_b_46_54536 = seg_13_17_sp4_r_v_b_11_54536;
  assign seg_14_14_sp4_v_b_47_54537 = seg_14_17_sp4_v_b_10_54537;
  assign seg_14_14_sp4_v_b_4_54162 = seg_13_13_sp4_r_v_b_17_54162;
  assign seg_14_14_sp4_v_b_5_54161 = seg_14_11_sp4_v_b_40_54161;
  assign seg_14_14_sp4_v_b_8_54166 = net_54166;
  assign seg_14_15_lutff_0_out_54502 = net_54502;
  assign seg_14_15_lutff_2_out_54504 = net_54504;
  assign seg_14_15_lutff_4_out_54506 = net_54506;
  assign seg_14_15_lutff_6_out_54508 = net_54508;
  assign seg_14_15_lutff_7_out_54509 = net_54509;
  assign seg_14_15_neigh_op_tnl_1_50795 = seg_13_16_lutff_1_out_50795;
  assign seg_14_15_sp4_h_r_14_54642 = net_54642;
  assign seg_14_15_sp4_r_v_b_23_58244 = net_58244;
  assign seg_14_15_sp4_v_b_0_54281 = seg_13_14_sp4_r_v_b_13_54281;
  assign seg_14_15_sp4_v_b_10_54291 = net_54291;
  assign seg_14_15_sp4_v_b_2_54283 = net_54283;
  assign seg_14_15_sp4_v_b_39_54652 = seg_13_17_sp4_r_v_b_15_54652;
  assign seg_14_15_sp4_v_b_3_54282 = seg_14_14_sp4_v_b_14_54282;
  assign seg_14_15_sp4_v_b_4_54285 = net_54285;
  assign seg_14_15_sp4_v_b_9_54288 = seg_14_14_sp4_v_b_20_54288;
  assign seg_14_15_sp4_v_t_41_54777 = seg_13_16_sp4_r_v_b_41_54777;
  assign seg_14_16_lutff_0_out_54625 = net_54625;
  assign seg_14_16_lutff_3_out_54628 = net_54628;
  assign seg_14_16_lutff_5_out_54630 = net_54630;
  assign seg_14_16_lutff_6_out_54631 = net_54631;
  assign seg_14_16_lutff_7_out_54632 = net_54632;
  assign seg_14_16_neigh_op_bot_0_54502 = seg_14_15_lutff_0_out_54502;
  assign seg_14_16_neigh_op_bot_4_54506 = seg_14_15_lutff_4_out_54506;
  assign seg_14_16_neigh_op_bot_7_54509 = seg_14_15_lutff_7_out_54509;
  assign seg_14_16_neigh_op_tnl_6_50923 = seg_13_17_lutff_6_out_50923;
  assign seg_14_16_sp4_h_r_32_50939 = seg_12_16_sp4_h_r_8_50939;
  assign seg_14_16_sp4_r_v_b_43_58609 = seg_15_19_sp4_v_b_6_58609;
  assign seg_14_16_sp4_v_b_2_54406 = net_54406;
  assign seg_14_16_sp4_v_b_8_54412 = net_54412;
  assign seg_14_16_sp4_v_t_41_54900 = seg_13_17_sp4_r_v_b_41_54900;
  assign seg_14_17_lutff_1_out_54749 = net_54749;
  assign seg_14_17_lutff_2_out_54750 = net_54750;
  assign seg_14_17_lutff_3_out_54751 = net_54751;
  assign seg_14_17_lutff_7_out_54755 = net_54755;
  assign seg_14_17_neigh_op_rgt_2_58580 = seg_15_17_lutff_2_out_58580;
  assign seg_14_17_neigh_op_rgt_7_58585 = seg_15_17_lutff_7_out_58585;
  assign seg_14_17_sp4_h_l_42_43399 = seg_11_17_sp4_h_r_18_43399;
  assign seg_14_17_sp4_h_l_43_43398 = seg_10_17_sp4_h_r_6_43398;
  assign seg_14_17_sp4_h_l_45_43400 = seg_10_17_sp4_h_r_8_43400;
  assign seg_14_17_sp4_r_v_b_30_58609 = seg_15_19_sp4_v_b_6_58609;
  assign seg_14_17_sp4_v_b_10_54537 = net_54537;
  assign seg_14_17_sp4_v_t_36_55018 = seg_13_19_sp4_r_v_b_25_55018;
  assign seg_14_18_lutff_0_out_54871 = net_54871;
  assign seg_14_18_lutff_1_out_54872 = net_54872;
  assign seg_14_18_lutff_3_out_54874 = net_54874;
  assign seg_14_18_lutff_5_out_54876 = net_54876;
  assign seg_14_18_neigh_op_lft_3_51043 = seg_13_18_lutff_3_out_51043;
  assign seg_14_18_neigh_op_lft_5_51045 = seg_13_18_lutff_5_out_51045;
  assign seg_14_18_neigh_op_tnr_3_58827 = seg_15_19_lutff_3_out_58827;
  assign seg_14_18_sp4_h_l_41_43519 = seg_10_18_sp4_h_r_4_43519;
  assign seg_14_18_sp4_h_l_45_43523 = seg_10_18_sp4_h_r_8_43523;
  assign seg_14_18_sp4_h_r_14_55011 = net_55011;
  assign seg_14_18_sp4_h_r_41_47350 = seg_11_18_sp4_h_r_4_47350;
  assign seg_14_18_sp4_h_r_8_58846 = net_58846;
  assign seg_14_18_sp4_h_r_9_58847 = seg_17_18_sp4_h_r_44_58847;
  assign seg_14_18_sp4_r_v_b_41_58853 = net_58853;
  assign seg_14_18_sp4_v_b_38_55020 = seg_14_20_sp4_v_b_14_55020;
  assign seg_14_19_lutff_0_out_54994 = net_54994;
  assign seg_14_19_lutff_1_out_54995 = net_54995;
  assign seg_14_19_lutff_6_out_55000 = net_55000;
  assign seg_14_19_lutff_7_out_55001 = net_55001;
  assign seg_14_19_neigh_op_rgt_3_58827 = seg_15_19_lutff_3_out_58827;
  assign seg_14_19_neigh_op_top_0_55117 = seg_14_20_lutff_0_out_55117;
  assign seg_14_19_neigh_op_top_4_55121 = seg_14_20_lutff_4_out_55121;
  assign seg_14_19_sp4_h_l_37_43636 = seg_10_19_sp4_h_r_0_43636;
  assign seg_14_19_sp4_h_l_39_43640 = seg_10_19_sp4_h_r_2_43640;
  assign seg_14_19_sp4_h_l_43_43644 = seg_10_19_sp4_h_r_6_43644;
  assign seg_14_19_sp4_h_l_47_43638 = seg_10_19_sp4_h_r_10_43638;
  assign seg_14_19_sp4_h_r_11_58962 = seg_15_19_sp4_h_r_22_58962;
  assign seg_14_19_sp4_h_r_43_47475 = seg_11_19_sp4_h_r_6_47475;
  assign seg_14_20_lutff_0_out_55117 = net_55117;
  assign seg_14_20_lutff_1_out_55118 = net_55118;
  assign seg_14_20_lutff_2_out_55119 = net_55119;
  assign seg_14_20_lutff_4_out_55121 = net_55121;
  assign seg_14_20_neigh_op_bnr_3_58827 = seg_15_19_lutff_3_out_58827;
  assign seg_14_20_neigh_op_lft_4_51290 = seg_13_20_lutff_4_out_51290;
  assign seg_14_20_neigh_op_lft_6_51292 = seg_13_20_lutff_6_out_51292;
  assign seg_14_20_neigh_op_top_7_55247 = seg_14_21_lutff_7_out_55247;
  assign seg_14_20_sp4_h_l_37_43759 = seg_10_20_sp4_h_r_0_43759;
  assign seg_14_20_sp4_h_l_39_43763 = seg_10_20_sp4_h_r_2_43763;
  assign seg_14_20_sp4_h_l_41_43765 = seg_10_20_sp4_h_r_4_43765;
  assign seg_14_20_sp4_h_l_43_43767 = seg_10_20_sp4_h_r_6_43767;
  assign seg_14_20_sp4_h_r_10_59084 = net_59084;
  assign seg_14_20_sp4_r_v_b_27_58973 = net_58973;
  assign seg_14_20_sp4_v_b_14_55020 = net_55020;
  assign seg_14_21_lutff_7_out_55247 = net_55247;
  assign seg_14_21_sp4_h_l_45_43892 = seg_12_21_sp4_h_r_32_43892;
  assign seg_14_21_sp4_h_r_1_59206 = seg_15_21_sp4_h_r_12_59206;
  assign seg_14_23_sp4_h_l_45_44138 = seg_12_23_sp4_h_r_32_44138;
  assign seg_14_26_lutff_3_out_55858 = net_55858;
  assign seg_14_26_sp4_r_v_b_25_59709 = net_59709;
  assign seg_14_27_lutff_2_out_55980 = net_55980;
  assign seg_14_27_lutff_5_out_55983 = net_55983;
  assign seg_14_27_neigh_op_lft_5_52152 = seg_13_27_lutff_5_out_52152;
  assign seg_14_27_sp4_h_r_36_48452 = seg_12_27_sp4_h_r_12_48452;
  assign seg_14_27_sp4_h_r_38_48456 = seg_12_27_sp4_h_r_14_48456;
  assign seg_14_27_sp4_r_v_b_10_59597 = seg_15_27_sp4_v_b_10_59597;
  assign seg_14_27_sp4_r_v_b_35_59842 = net_59842;
  assign seg_14_28_neigh_op_rgt_0_59931 = seg_15_28_lutff_0_out_59931;
  assign seg_14_28_sp4_h_r_18_56245 = net_56245;
  assign seg_14_28_sp4_h_r_34_52407 = net_52407;
  assign seg_14_28_sp4_v_b_0_55880 = seg_13_27_sp4_r_v_b_13_55880;
  assign seg_14_2_lutff_2_out_52869 = net_52869;
  assign seg_14_2_lutff_3_out_52870 = net_52870;
  assign seg_14_2_neigh_op_rgt_0_56697 = seg_15_2_lutff_0_out_56697;
  assign seg_14_2_neigh_op_tnr_2_56858 = seg_15_3_lutff_2_out_56858;
  assign seg_14_2_neigh_op_tnr_3_56859 = seg_15_3_lutff_3_out_56859;
  assign seg_14_2_neigh_op_tnr_7_56863 = seg_15_3_lutff_7_out_56863;
  assign seg_14_2_neigh_op_top_3_53029 = seg_14_3_lutff_3_out_53029;
  assign seg_14_2_sp12_v_b_12_56584 = net_56584;
  assign seg_14_2_sp4_h_r_10_56870 = net_56870;
  assign seg_14_3_lutff_0_out_53026 = net_53026;
  assign seg_14_3_lutff_1_out_53027 = net_53027;
  assign seg_14_3_lutff_2_out_53028 = net_53028;
  assign seg_14_3_lutff_3_out_53029 = net_53029;
  assign seg_14_3_lutff_4_out_53030 = net_53030;
  assign seg_14_3_lutff_5_out_53031 = net_53031;
  assign seg_14_3_lutff_6_out_53032 = net_53032;
  assign seg_14_3_lutff_7_out_53033 = net_53033;
  assign seg_14_3_neigh_op_bnr_0_56697 = seg_15_2_lutff_0_out_56697;
  assign seg_14_3_neigh_op_bnr_1_56698 = seg_15_2_lutff_1_out_56698;
  assign seg_14_3_neigh_op_lft_7_49202 = seg_13_3_lutff_7_out_49202;
  assign seg_14_3_neigh_op_rgt_2_56858 = seg_15_3_lutff_2_out_56858;
  assign seg_14_3_neigh_op_rgt_3_56859 = seg_15_3_lutff_3_out_56859;
  assign seg_14_3_neigh_op_rgt_7_56863 = seg_15_3_lutff_7_out_56863;
  assign seg_14_3_neigh_op_top_0_53149 = seg_14_4_lutff_0_out_53149;
  assign seg_14_3_neigh_op_top_1_53150 = seg_14_4_lutff_1_out_53150;
  assign seg_14_3_neigh_op_top_4_53153 = seg_14_4_lutff_4_out_53153;
  assign seg_14_3_neigh_op_top_7_53156 = seg_14_4_lutff_7_out_53156;
  assign seg_14_3_sp12_v_b_11_56584 = seg_14_2_sp12_v_b_12_56584;
  assign seg_14_3_sp4_v_b_19_52929 = seg_13_3_sp4_r_v_b_19_52929;
  assign seg_14_4_lutff_0_out_53149 = net_53149;
  assign seg_14_4_lutff_1_out_53150 = net_53150;
  assign seg_14_4_lutff_2_out_53151 = net_53151;
  assign seg_14_4_lutff_4_out_53153 = net_53153;
  assign seg_14_4_lutff_5_out_53154 = net_53154;
  assign seg_14_4_lutff_7_out_53156 = net_53156;
  assign seg_14_4_neigh_op_bot_0_53026 = seg_14_3_lutff_0_out_53026;
  assign seg_14_4_neigh_op_bot_6_53032 = seg_14_3_lutff_6_out_53032;
  assign seg_14_4_neigh_op_lft_2_49320 = seg_13_4_lutff_2_out_49320;
  assign seg_14_4_neigh_op_lft_3_49321 = seg_13_4_lutff_3_out_49321;
  assign seg_14_7_lutff_1_out_53519 = net_53519;
  assign seg_14_7_lutff_6_out_53524 = net_53524;
  assign seg_14_7_lutff_7_out_53525 = net_53525;
  assign seg_14_7_sp4_h_l_47_42162 = seg_10_7_sp4_h_r_10_42162;
  assign seg_14_7_sp4_v_b_28_53547 = net_53547;
  assign seg_14_8_lutff_6_out_53647 = net_53647;
  assign seg_14_8_lutff_7_out_53648 = net_53648;
  assign seg_14_8_neigh_op_bot_6_53524 = seg_14_7_lutff_6_out_53524;
  assign seg_14_8_neigh_op_lft_3_49813 = seg_13_8_lutff_3_out_49813;
  assign seg_14_8_neigh_op_tnl_0_49933 = seg_13_9_lutff_0_out_49933;
  assign seg_14_8_neigh_op_tnl_5_49938 = seg_13_9_lutff_5_out_49938;
  assign seg_14_8_neigh_op_top_3_53767 = seg_14_9_lutff_3_out_53767;
  assign seg_14_8_neigh_op_top_6_53770 = seg_14_9_lutff_6_out_53770;
  assign seg_14_8_sp4_h_r_25_49946 = seg_13_8_sp4_h_r_12_49946;
  assign seg_14_8_sp4_h_r_8_57616 = net_57616;
  assign seg_14_8_sp4_r_v_b_11_57259 = net_57259;
  assign seg_14_8_sp4_r_v_b_25_57495 = net_57495;
  assign seg_14_9_lutff_2_out_53766 = net_53766;
  assign seg_14_9_lutff_3_out_53767 = net_53767;
  assign seg_14_9_lutff_4_out_53768 = net_53768;
  assign seg_14_9_lutff_5_out_53769 = net_53769;
  assign seg_14_9_lutff_6_out_53770 = net_53770;
  assign seg_14_9_lutff_7_out_53771 = net_53771;
  assign seg_14_9_neigh_op_bnr_0_57471 = seg_15_8_lutff_0_out_57471;
  assign seg_14_9_neigh_op_bot_6_53647 = seg_14_8_lutff_6_out_53647;
  assign seg_14_9_neigh_op_bot_7_53648 = seg_14_8_lutff_7_out_53648;
  assign seg_14_9_neigh_op_lft_0_49933 = seg_13_9_lutff_0_out_49933;
  assign seg_14_9_neigh_op_lft_1_49934 = seg_13_9_lutff_1_out_49934;
  assign seg_14_9_neigh_op_lft_5_49938 = seg_13_9_lutff_5_out_49938;
  assign seg_14_9_neigh_op_lft_6_49939 = seg_13_9_lutff_6_out_49939;
  assign seg_14_9_sp4_v_b_4_53547 = seg_14_7_sp4_v_b_28_53547;
  assign seg_15_0_span4_vert_19_56732 = seg_15_2_sp4_v_b_6_56732;
  assign seg_15_10_lutff_4_out_57721 = net_57721;
  assign seg_15_10_neigh_op_bnr_6_61430 = seg_16_9_lutff_6_out_61430;
  assign seg_15_10_neigh_op_bot_0_57594 = seg_15_9_lutff_0_out_57594;
  assign seg_15_10_neigh_op_bot_5_57599 = seg_15_9_lutff_5_out_57599;
  assign seg_15_10_neigh_op_rgt_5_61552 = seg_16_10_lutff_5_out_61552;
  assign seg_15_10_sp12_v_b_12_60943 = net_60943;
  assign seg_15_10_sp12_v_b_20_61435 = seg_15_20_sp12_v_b_0_61435;
  assign seg_15_10_sp4_h_l_45_46370 = seg_11_10_sp4_h_r_8_46370;
  assign seg_15_10_sp4_h_r_20_57863 = net_57863;
  assign seg_15_10_sp4_h_r_24_54022 = net_54022;
  assign seg_15_10_sp4_h_r_3_61687 = seg_18_10_sp4_h_r_38_61687;
  assign seg_15_10_sp4_h_r_8_61692 = net_61692;
  assign seg_15_10_sp4_r_v_b_41_61699 = net_61699;
  assign seg_15_10_sp4_r_v_b_9_61333 = net_61333;
  assign seg_15_10_sp4_v_b_19_57625 = seg_15_9_sp4_v_b_30_57625;
  assign seg_15_10_sp4_v_b_1_57495 = seg_14_8_sp4_r_v_b_25_57495;
  assign seg_15_10_sp4_v_b_24_57742 = net_57742;
  assign seg_15_10_sp4_v_b_40_57868 = net_57868;
  assign seg_15_10_sp4_v_b_42_57870 = net_57870;
  assign seg_15_11_lutff_1_out_57841 = net_57841;
  assign seg_15_11_lutff_2_out_57842 = net_57842;
  assign seg_15_11_lutff_4_out_57844 = net_57844;
  assign seg_15_11_lutff_6_out_57846 = net_57846;
  assign seg_15_11_lutff_7_out_57847 = net_57847;
  assign seg_15_11_neigh_op_bnr_5_61552 = seg_16_10_lutff_5_out_61552;
  assign seg_15_11_neigh_op_lft_0_54010 = seg_14_11_lutff_0_out_54010;
  assign seg_15_11_neigh_op_lft_5_54015 = seg_14_11_lutff_5_out_54015;
  assign seg_15_11_neigh_op_lft_6_54016 = seg_14_11_lutff_6_out_54016;
  assign seg_15_11_neigh_op_rgt_0_61670 = seg_16_11_lutff_0_out_61670;
  assign seg_15_11_neigh_op_rgt_1_61671 = seg_16_11_lutff_1_out_61671;
  assign seg_15_11_neigh_op_rgt_4_61674 = seg_16_11_lutff_4_out_61674;
  assign seg_15_11_sp12_v_b_10_60942 = seg_15_9_sp12_v_b_14_60942;
  assign seg_15_11_sp4_h_r_22_57978 = net_57978;
  assign seg_15_11_sp4_r_v_b_20_61579 = seg_16_9_sp4_v_b_44_61579;
  assign seg_15_11_sp4_r_v_b_27_61696 = net_61696;
  assign seg_15_12_lutff_0_out_57963 = net_57963;
  assign seg_15_12_lutff_1_out_57964 = net_57964;
  assign seg_15_12_lutff_2_out_57965 = net_57965;
  assign seg_15_12_lutff_3_out_57966 = net_57966;
  assign seg_15_12_lutff_4_out_57967 = net_57967;
  assign seg_15_12_lutff_5_out_57968 = net_57968;
  assign seg_15_12_lutff_6_out_57969 = net_57969;
  assign seg_15_12_lutff_7_out_57970 = net_57970;
  assign seg_15_12_neigh_op_top_3_58089 = seg_15_13_lutff_3_out_58089;
  assign seg_15_12_neigh_op_top_4_58090 = seg_15_13_lutff_4_out_58090;
  assign seg_15_12_sp4_h_l_41_46612 = seg_13_12_sp4_h_r_28_46612;
  assign seg_15_12_sp4_h_l_45_46616 = seg_11_12_sp4_h_r_8_46616;
  assign seg_15_12_sp4_r_v_b_31_61823 = seg_15_14_sp4_r_v_b_7_61823;
  assign seg_15_12_sp4_v_b_0_57742 = seg_15_10_sp4_v_b_24_57742;
  assign seg_15_12_sp4_v_b_11_57751 = seg_15_9_sp4_v_b_46_57751;
  assign seg_15_12_sp4_v_b_28_57992 = seg_15_14_sp4_v_b_4_57992;
  assign seg_15_12_sp4_v_b_36_58110 = seg_15_14_sp4_v_b_12_58110;
  assign seg_15_12_sp4_v_b_47_58121 = seg_14_14_sp4_r_v_b_23_58121;
  assign seg_15_12_sp4_v_t_46_58243 = seg_15_15_sp4_v_b_22_58243;
  assign seg_15_12_sp4_v_t_47_58244 = seg_14_15_sp4_r_v_b_23_58244;
  assign seg_15_13_lutff_3_out_58089 = net_58089;
  assign seg_15_13_lutff_4_out_58090 = net_58090;
  assign seg_15_13_lutff_7_out_58093 = net_58093;
  assign seg_15_13_neigh_op_bot_0_57963 = seg_15_12_lutff_0_out_57963;
  assign seg_15_13_neigh_op_bot_2_57965 = seg_15_12_lutff_2_out_57965;
  assign seg_15_13_neigh_op_bot_4_57967 = seg_15_12_lutff_4_out_57967;
  assign seg_15_13_neigh_op_bot_5_57968 = seg_15_12_lutff_5_out_57968;
  assign seg_15_13_neigh_op_tnl_1_54380 = seg_14_14_lutff_1_out_54380;
  assign seg_15_13_neigh_op_top_0_58209 = seg_15_14_lutff_0_out_58209;
  assign seg_15_13_neigh_op_top_5_58214 = seg_15_14_lutff_5_out_58214;
  assign seg_15_13_sp4_h_l_43_46737 = seg_13_13_sp4_h_r_30_46737;
  assign seg_15_13_sp4_h_r_0_62051 = net_62051;
  assign seg_15_13_sp4_h_r_10_62053 = net_62053;
  assign seg_15_13_sp4_h_r_12_58222 = net_58222;
  assign seg_15_13_sp4_h_r_18_58230 = net_58230;
  assign seg_15_13_sp4_h_r_28_54397 = seg_13_13_sp4_h_r_4_54397;
  assign seg_15_13_sp4_h_r_4_62057 = net_62057;
  assign seg_15_13_sp4_r_v_b_13_61818 = net_61818;
  assign seg_15_13_sp4_r_v_b_19_61824 = net_61824;
  assign seg_15_13_sp4_r_v_b_3_61696 = seg_15_11_sp4_r_v_b_27_61696;
  assign seg_15_13_sp4_r_v_b_4_61699 = seg_15_10_sp4_r_v_b_41_61699;
  assign seg_15_13_sp4_v_b_2_57867 = seg_14_12_sp4_r_v_b_15_57867;
  assign seg_15_13_sp4_v_b_37_58234 = seg_15_16_sp4_v_b_0_58234;
  assign seg_15_13_sp4_v_b_43_58240 = seg_15_16_sp4_v_b_6_58240;
  assign seg_15_13_sp4_v_t_38_58358 = seg_15_16_sp4_v_b_14_58358;
  assign seg_15_14_lutff_0_out_58209 = net_58209;
  assign seg_15_14_lutff_5_out_58214 = net_58214;
  assign seg_15_14_neigh_op_bnl_2_54258 = seg_14_13_lutff_2_out_54258;
  assign seg_15_14_neigh_op_lft_6_54385 = seg_14_14_lutff_6_out_54385;
  assign seg_15_14_neigh_op_top_1_58333 = seg_15_15_lutff_1_out_58333;
  assign seg_15_14_neigh_op_top_7_58339 = seg_15_15_lutff_7_out_58339;
  assign seg_15_14_sp12_v_b_4_60943 = seg_15_10_sp12_v_b_12_60943;
  assign seg_15_14_sp4_h_l_38_46857 = seg_12_14_sp4_h_r_14_46857;
  assign seg_15_14_sp4_h_r_14_58349 = net_58349;
  assign seg_15_14_sp4_h_r_2_62178 = net_62178;
  assign seg_15_14_sp4_h_r_41_50689 = seg_12_14_sp4_h_r_4_50689;
  assign seg_15_14_sp4_h_r_8_62184 = net_62184;
  assign seg_15_14_sp4_r_v_b_15_61943 = net_61943;
  assign seg_15_14_sp4_r_v_b_19_61947 = net_61947;
  assign seg_15_14_sp4_r_v_b_33_62071 = seg_15_16_sp4_r_v_b_9_62071;
  assign seg_15_14_sp4_r_v_b_7_61823 = net_61823;
  assign seg_15_14_sp4_v_b_0_57988 = seg_14_11_sp4_r_v_b_37_57988;
  assign seg_15_14_sp4_v_b_12_58110 = net_58110;
  assign seg_15_14_sp4_v_b_47_58367 = seg_15_17_sp4_v_b_10_58367;
  assign seg_15_14_sp4_v_b_4_57992 = net_57992;
  assign seg_15_14_sp4_v_b_7_57993 = seg_14_12_sp4_r_v_b_31_57993;
  assign seg_15_14_sp4_v_b_9_57995 = seg_14_12_sp4_r_v_b_33_57995;
  assign seg_15_14_sp4_v_t_46_58489 = seg_15_17_sp4_v_b_22_58489;
  assign seg_15_15_lutff_0_out_58332 = net_58332;
  assign seg_15_15_lutff_1_out_58333 = net_58333;
  assign seg_15_15_lutff_5_out_58337 = net_58337;
  assign seg_15_15_lutff_7_out_58339 = net_58339;
  assign seg_15_15_neigh_op_tnl_5_54630 = seg_14_16_lutff_5_out_54630;
  assign seg_15_15_sp4_h_l_39_46979 = seg_13_15_sp4_h_r_26_46979;
  assign seg_15_15_sp4_h_r_26_54641 = seg_13_15_sp4_h_r_2_54641;
  assign seg_15_15_sp4_h_r_41_50812 = seg_12_15_sp4_h_r_4_50812;
  assign seg_15_15_sp4_h_r_4_62303 = net_62303;
  assign seg_15_15_sp4_h_r_8_62307 = net_62307;
  assign seg_15_15_sp4_r_v_b_13_62064 = net_62064;
  assign seg_15_15_sp4_v_b_22_58243 = net_58243;
  assign seg_15_15_sp4_v_b_26_58359 = seg_15_17_sp4_v_b_2_58359;
  assign seg_15_15_sp4_v_t_43_58609 = seg_15_19_sp4_v_b_6_58609;
  assign seg_15_16_lutff_6_out_58461 = net_58461;
  assign seg_15_16_neigh_op_rgt_2_62287 = seg_16_16_lutff_2_out_62287;
  assign seg_15_16_sp4_h_l_39_47102 = seg_13_16_sp4_h_r_26_47102;
  assign seg_15_16_sp4_h_r_26_54764 = net_54764;
  assign seg_15_16_sp4_h_r_6_62428 = seg_17_16_sp4_h_r_30_62428;
  assign seg_15_16_sp4_r_v_b_9_62071 = net_62071;
  assign seg_15_16_sp4_v_b_0_58234 = net_58234;
  assign seg_15_16_sp4_v_b_14_58358 = net_58358;
  assign seg_15_16_sp4_v_b_2_58236 = seg_14_13_sp4_r_v_b_39_58236;
  assign seg_15_16_sp4_v_b_43_58609 = seg_15_19_sp4_v_b_6_58609;
  assign seg_15_16_sp4_v_b_6_58240 = net_58240;
  assign seg_15_16_sp4_v_b_9_58241 = seg_14_14_sp4_r_v_b_33_58241;
  assign seg_15_16_sp4_v_t_37_58726 = seg_15_20_sp4_v_b_0_58726;
  assign seg_15_16_sp4_v_t_46_58735 = seg_15_19_sp4_v_b_22_58735;
  assign seg_15_17_lutff_0_out_58578 = net_58578;
  assign seg_15_17_lutff_2_out_58580 = net_58580;
  assign seg_15_17_lutff_7_out_58585 = net_58585;
  assign seg_15_17_sp4_h_r_28_54889 = net_54889;
  assign seg_15_17_sp4_v_b_10_58367 = net_58367;
  assign seg_15_17_sp4_v_b_22_58489 = net_58489;
  assign seg_15_17_sp4_v_b_2_58359 = net_58359;
  assign seg_15_17_sp4_v_b_30_58609 = seg_15_19_sp4_v_b_6_58609;
  assign seg_15_17_sp4_v_b_37_58726 = seg_15_20_sp4_v_b_0_58726;
  assign seg_15_17_sp4_v_t_38_58850 = seg_15_20_sp4_v_b_14_58850;
  assign seg_15_17_sp4_v_t_40_58852 = seg_15_20_sp4_v_b_16_58852;
  assign seg_15_17_sp4_v_t_41_58853 = seg_14_18_sp4_r_v_b_41_58853;
  assign seg_15_18_lutff_1_out_58702 = net_58702;
  assign seg_15_18_lutff_2_out_58703 = net_58703;
  assign seg_15_18_lutff_4_out_58705 = net_58705;
  assign seg_15_18_lutff_7_out_58708 = net_58708;
  assign seg_15_18_neigh_op_tnl_1_54995 = seg_14_19_lutff_1_out_54995;
  assign seg_15_18_neigh_op_top_0_58824 = seg_15_19_lutff_0_out_58824;
  assign seg_15_18_neigh_op_top_6_58830 = seg_15_19_lutff_6_out_58830;
  assign seg_15_18_sp12_h_r_0_62662 = seg_17_18_sp12_h_r_4_62662;
  assign seg_15_18_sp4_h_l_39_47348 = seg_11_18_sp4_h_r_2_47348;
  assign seg_15_18_sp4_h_l_40_47351 = seg_12_18_sp4_h_r_16_47351;
  assign seg_15_18_sp4_h_r_0_62666 = net_62666;
  assign seg_15_18_sp4_h_r_12_58837 = net_58837;
  assign seg_15_18_sp4_v_b_24_58726 = seg_15_20_sp4_v_b_0_58726;
  assign seg_15_18_sp4_v_t_36_58971 = seg_15_21_sp4_v_b_12_58971;
  assign seg_15_18_sp4_v_t_38_58973 = seg_14_20_sp4_r_v_b_27_58973;
  assign seg_15_18_sp4_v_t_45_58980 = seg_15_22_sp4_v_b_8_58980;
  assign seg_15_19_lutff_0_out_58824 = net_58824;
  assign seg_15_19_lutff_3_out_58827 = net_58827;
  assign seg_15_19_lutff_5_out_58829 = net_58829;
  assign seg_15_19_lutff_6_out_58830 = net_58830;
  assign seg_15_19_neigh_op_top_0_58947 = seg_15_20_lutff_0_out_58947;
  assign seg_15_19_sp4_h_r_22_58962 = net_58962;
  assign seg_15_19_sp4_h_r_38_51303 = net_51303;
  assign seg_15_19_sp4_h_r_6_62797 = net_62797;
  assign seg_15_19_sp4_r_v_b_23_62566 = net_62566;
  assign seg_15_19_sp4_r_v_b_7_62438 = net_62438;
  assign seg_15_19_sp4_v_b_22_58735 = net_58735;
  assign seg_15_19_sp4_v_b_6_58609 = net_58609;
  assign seg_15_20_lutff_0_out_58947 = net_58947;
  assign seg_15_20_lutff_2_out_58949 = net_58949;
  assign seg_15_20_neigh_op_bot_3_58827 = seg_15_19_lutff_3_out_58827;
  assign seg_15_20_sp12_v_b_0_61435 = net_61435;
  assign seg_15_20_sp4_h_r_30_55260 = net_55260;
  assign seg_15_20_sp4_h_r_44_51432 = net_51432;
  assign seg_15_20_sp4_r_v_b_1_62555 = net_62555;
  assign seg_15_20_sp4_v_b_0_58726 = net_58726;
  assign seg_15_20_sp4_v_b_14_58850 = net_58850;
  assign seg_15_20_sp4_v_b_16_58852 = net_58852;
  assign seg_15_20_sp4_v_b_47_59105 = seg_15_23_sp4_v_b_10_59105;
  assign seg_15_20_sp4_v_t_37_59218 = seg_15_22_sp4_v_b_24_59218;
  assign seg_15_20_sp4_v_t_38_59219 = seg_15_23_sp4_v_b_14_59219;
  assign seg_15_21_sp4_h_l_38_47718 = seg_12_21_sp4_h_r_14_47718;
  assign seg_15_21_sp4_h_l_44_47724 = seg_12_21_sp4_h_r_20_47724;
  assign seg_15_21_sp4_h_r_12_59206 = net_59206;
  assign seg_15_21_sp4_h_r_28_55381 = net_55381;
  assign seg_15_21_sp4_h_r_44_51555 = net_51555;
  assign seg_15_21_sp4_r_v_b_13_62802 = net_62802;
  assign seg_15_21_sp4_v_b_12_58971 = net_58971;
  assign seg_15_21_sp4_v_b_34_59105 = seg_15_23_sp4_v_b_10_59105;
  assign seg_15_22_lutff_4_out_59197 = net_59197;
  assign seg_15_22_lutff_5_out_59198 = net_59198;
  assign seg_15_22_sp4_v_b_24_59218 = net_59218;
  assign seg_15_22_sp4_v_b_8_58980 = net_58980;
  assign seg_15_23_lutff_1_out_59317 = net_59317;
  assign seg_15_23_neigh_op_bot_5_59198 = seg_15_22_lutff_5_out_59198;
  assign seg_15_23_sp4_h_r_42_51799 = net_51799;
  assign seg_15_23_sp4_v_b_10_59105 = net_59105;
  assign seg_15_23_sp4_v_b_14_59219 = net_59219;
  assign seg_15_23_sp4_v_b_34_59351 = seg_15_25_sp4_v_b_10_59351;
  assign seg_15_23_sp4_v_t_39_59589 = seg_15_25_sp4_v_b_26_59589;
  assign seg_15_25_sp4_r_v_b_11_63180 = net_63180;
  assign seg_15_25_sp4_r_v_b_27_63418 = net_63418;
  assign seg_15_25_sp4_v_b_10_59351 = net_59351;
  assign seg_15_25_sp4_v_b_26_59589 = net_59589;
  assign seg_15_25_sp4_v_t_42_59838 = seg_15_28_sp4_v_b_18_59838;
  assign seg_15_27_neigh_op_top_4_59935 = seg_15_28_lutff_4_out_59935;
  assign seg_15_27_sp4_v_b_10_59597 = net_59597;
  assign seg_15_28_lutff_0_out_59931 = net_59931;
  assign seg_15_28_lutff_4_out_59935 = net_59935;
  assign seg_15_28_lutff_5_out_59936 = net_59936;
  assign seg_15_28_neigh_op_rgt_1_63762 = seg_16_28_lutff_1_out_63762;
  assign seg_15_28_neigh_op_rgt_3_63764 = seg_16_28_lutff_3_out_63764;
  assign seg_15_28_neigh_op_rgt_5_63766 = seg_16_28_lutff_5_out_63766;
  assign seg_15_28_neigh_op_rgt_6_63767 = seg_16_28_lutff_6_out_63767;
  assign seg_15_28_sp4_h_l_42_48583 = seg_12_28_sp4_h_r_18_48583;
  assign seg_15_28_sp4_h_r_30_56244 = net_56244;
  assign seg_15_28_sp4_h_r_46_52408 = net_52408;
  assign seg_15_28_sp4_v_b_18_59838 = net_59838;
  assign seg_15_28_sp4_v_b_1_59709 = seg_14_26_sp4_r_v_b_25_59709;
  assign seg_15_29_lutff_5_out_60059 = net_60059;
  assign seg_15_29_neigh_op_bnr_1_63762 = seg_16_28_lutff_1_out_63762;
  assign seg_15_29_neigh_op_bnr_3_63764 = seg_16_28_lutff_3_out_63764;
  assign seg_15_29_neigh_op_bnr_5_63766 = seg_16_28_lutff_5_out_63766;
  assign seg_15_29_neigh_op_bnr_6_63767 = seg_16_28_lutff_6_out_63767;
  assign seg_15_29_sp4_r_v_b_31_63914 = net_63914;
  assign seg_15_29_sp4_v_b_11_59842 = seg_14_27_sp4_r_v_b_35_59842;
  assign seg_15_2_lutff_0_out_56697 = net_56697;
  assign seg_15_2_lutff_1_out_56698 = net_56698;
  assign seg_15_2_lutff_2_out_56699 = net_56699;
  assign seg_15_2_lutff_6_out_56703 = net_56703;
  assign seg_15_2_neigh_op_top_2_56858 = seg_15_3_lutff_2_out_56858;
  assign seg_15_2_neigh_op_top_3_56859 = seg_15_3_lutff_3_out_56859;
  assign seg_15_2_neigh_op_top_7_56863 = seg_15_3_lutff_7_out_56863;
  assign seg_15_2_sp4_v_b_6_56732 = net_56732;
  assign seg_15_30_sp4_h_l_43_48824 = seg_11_30_sp4_h_r_6_48824;
  assign seg_15_3_lutff_1_out_56857 = net_56857;
  assign seg_15_3_lutff_2_out_56858 = net_56858;
  assign seg_15_3_lutff_3_out_56859 = net_56859;
  assign seg_15_3_lutff_4_out_56860 = net_56860;
  assign seg_15_3_lutff_6_out_56862 = net_56862;
  assign seg_15_3_lutff_7_out_56863 = net_56863;
  assign seg_15_3_neigh_op_bnr_5_60532 = seg_16_2_lutff_5_out_60532;
  assign seg_15_3_neigh_op_bot_0_56697 = seg_15_2_lutff_0_out_56697;
  assign seg_15_3_neigh_op_bot_2_56699 = seg_15_2_lutff_2_out_56699;
  assign seg_15_3_neigh_op_lft_4_53030 = seg_14_3_lutff_4_out_53030;
  assign seg_15_3_neigh_op_lft_5_53031 = seg_14_3_lutff_5_out_53031;
  assign seg_15_3_sp4_r_v_b_43_60840 = net_60840;
  assign seg_15_6_sp4_h_r_36_49700 = net_49700;
  assign seg_15_6_sp4_r_v_b_21_60965 = net_60965;
  assign seg_15_6_sp4_r_v_b_37_61203 = net_61203;
  assign seg_15_8_lutff_0_out_57471 = net_57471;
  assign seg_15_8_sp4_h_r_32_53786 = net_53786;
  assign seg_15_8_sp4_r_v_b_17_61207 = net_61207;
  assign seg_15_8_sp4_v_b_11_57259 = seg_14_8_sp4_r_v_b_11_57259;
  assign seg_15_9_lutff_0_out_57594 = net_57594;
  assign seg_15_9_lutff_5_out_57599 = net_57599;
  assign seg_15_9_neigh_op_rgt_2_61426 = seg_16_9_lutff_2_out_61426;
  assign seg_15_9_neigh_op_rgt_5_61429 = seg_16_9_lutff_5_out_61429;
  assign seg_15_9_sp12_v_b_14_60942 = net_60942;
  assign seg_15_9_sp12_v_b_23_61435 = seg_15_20_sp12_v_b_0_61435;
  assign seg_15_9_sp4_r_v_b_0_61203 = seg_15_6_sp4_r_v_b_37_61203;
  assign seg_15_9_sp4_r_v_b_36_61571 = seg_16_9_sp4_v_b_36_61571;
  assign seg_15_9_sp4_v_b_30_57625 = net_57625;
  assign seg_15_9_sp4_v_b_46_57751 = net_57751;
  assign seg_15_9_sp4_v_t_42_57870 = seg_15_10_sp4_v_b_42_57870;
  assign seg_16_10_lutff_5_out_61552 = net_61552;
  assign seg_16_10_neigh_op_bnr_1_65256 = seg_17_9_lutff_1_out_65256;
  assign seg_16_10_sp4_v_b_9_61333 = seg_15_10_sp4_r_v_b_9_61333;
  assign seg_16_11_lutff_0_out_61670 = net_61670;
  assign seg_16_11_lutff_1_out_61671 = net_61671;
  assign seg_16_11_lutff_4_out_61674 = net_61674;
  assign seg_16_11_lutff_5_out_61675 = net_61675;
  assign seg_16_11_neigh_op_top_2_61795 = seg_16_12_lutff_2_out_61795;
  assign seg_16_12_lutff_2_out_61795 = net_61795;
  assign seg_16_12_neigh_op_bnl_4_57844 = seg_15_11_lutff_4_out_57844;
  assign seg_16_12_neigh_op_bnl_6_57846 = seg_15_11_lutff_6_out_57846;
  assign seg_16_12_neigh_op_bot_5_61675 = seg_16_11_lutff_5_out_61675;
  assign seg_16_12_neigh_op_top_4_61920 = seg_16_13_lutff_4_out_61920;
  assign seg_16_12_sp4_h_r_0_65759 = net_65759;
  assign seg_16_12_sp4_h_r_12_61929 = net_61929;
  assign seg_16_12_sp4_h_r_26_58102 = seg_14_12_sp4_h_r_2_58102;
  assign seg_16_12_sp4_h_r_2_65763 = net_65763;
  assign seg_16_12_sp4_h_r_40_54275 = net_54275;
  assign seg_16_12_sp4_h_r_43_54276 = seg_13_12_sp4_h_r_6_54276;
  assign seg_16_12_sp4_r_v_b_35_65658 = net_65658;
  assign seg_16_12_sp4_v_b_17_61699 = seg_15_10_sp4_r_v_b_41_61699;
  assign seg_16_12_sp4_v_b_32_61826 = net_61826;
  assign seg_16_12_sp4_v_b_38_61942 = seg_16_14_sp4_v_b_14_61942;
  assign seg_16_12_sp4_v_b_42_61946 = net_61946;
  assign seg_16_12_sp4_v_b_45_61949 = seg_16_15_sp4_v_b_8_61949;
  assign seg_16_12_sp4_v_t_37_62064 = seg_15_15_sp4_r_v_b_13_62064;
  assign seg_16_12_sp4_v_t_39_62066 = seg_16_16_sp4_v_b_2_62066;
  assign seg_16_13_lutff_0_out_61916 = net_61916;
  assign seg_16_13_lutff_2_out_61918 = net_61918;
  assign seg_16_13_lutff_3_out_61919 = net_61919;
  assign seg_16_13_lutff_4_out_61920 = net_61920;
  assign seg_16_13_neigh_op_bnl_3_57966 = seg_15_12_lutff_3_out_57966;
  assign seg_16_13_neigh_op_top_5_62044 = seg_16_14_lutff_5_out_62044;
  assign seg_16_13_sp4_h_l_37_50560 = seg_14_13_sp4_h_r_24_50560;
  assign seg_16_13_sp4_h_l_39_50564 = seg_14_13_sp4_h_r_26_50564;
  assign seg_16_13_sp4_h_l_40_50567 = seg_13_13_sp4_h_r_16_50567;
  assign seg_16_13_sp4_h_r_26_58225 = seg_14_13_sp4_h_r_2_58225;
  assign seg_16_13_sp4_h_r_4_65888 = net_65888;
  assign seg_16_13_sp4_v_b_4_61699 = seg_15_10_sp4_r_v_b_41_61699;
  assign seg_16_14_lutff_1_out_62040 = net_62040;
  assign seg_16_14_lutff_5_out_62044 = net_62044;
  assign seg_16_14_lutff_7_out_62046 = net_62046;
  assign seg_16_14_sp4_v_b_0_61818 = seg_15_13_sp4_r_v_b_13_61818;
  assign seg_16_14_sp4_v_b_14_61942 = net_61942;
  assign seg_16_14_sp4_v_b_26_62066 = seg_16_16_sp4_v_b_2_62066;
  assign seg_16_14_sp4_v_b_6_61824 = seg_15_13_sp4_r_v_b_19_61824;
  assign seg_16_14_sp4_v_b_8_61826 = seg_16_12_sp4_v_b_32_61826;
  assign seg_16_14_sp4_v_t_47_62320 = seg_16_16_sp4_v_b_34_62320;
  assign seg_16_15_lutff_0_out_62162 = net_62162;
  assign seg_16_15_lutff_3_out_62165 = net_62165;
  assign seg_16_15_lutff_7_out_62169 = net_62169;
  assign seg_16_15_neigh_op_bot_1_62040 = seg_16_14_lutff_1_out_62040;
  assign seg_16_15_neigh_op_lft_7_58339 = seg_15_15_lutff_7_out_58339;
  assign seg_16_15_neigh_op_top_2_62287 = seg_16_16_lutff_2_out_62287;
  assign seg_16_15_sp4_h_l_38_50811 = seg_13_15_sp4_h_r_14_50811;
  assign seg_16_15_sp4_h_l_40_50813 = seg_13_15_sp4_h_r_16_50813;
  assign seg_16_15_sp4_h_r_10_66130 = net_66130;
  assign seg_16_15_sp4_h_r_12_62298 = net_62298;
  assign seg_16_15_sp4_h_r_38_54642 = seg_14_15_sp4_h_r_14_54642;
  assign seg_16_15_sp4_h_r_4_66134 = net_66134;
  assign seg_16_15_sp4_r_v_b_15_65897 = net_65897;
  assign seg_16_15_sp4_r_v_b_21_65903 = net_65903;
  assign seg_16_15_sp4_v_b_26_62189 = net_62189;
  assign seg_16_15_sp4_v_b_2_61943 = seg_15_14_sp4_r_v_b_15_61943;
  assign seg_16_15_sp4_v_b_6_61947 = seg_15_14_sp4_r_v_b_19_61947;
  assign seg_16_15_sp4_v_b_7_61946 = seg_16_12_sp4_v_b_42_61946;
  assign seg_16_15_sp4_v_b_8_61949 = net_61949;
  assign seg_16_15_sp4_v_t_42_62438 = seg_15_19_sp4_r_v_b_7_62438;
  assign seg_16_16_lutff_1_out_62286 = net_62286;
  assign seg_16_16_lutff_2_out_62287 = net_62287;
  assign seg_16_16_sp12_v_b_1_64773 = seg_16_9_sp12_v_b_14_64773;
  assign seg_16_16_sp4_h_r_2_66255 = net_66255;
  assign seg_16_16_sp4_h_r_3_66256 = seg_17_16_sp4_h_r_14_66256;
  assign seg_16_16_sp4_r_v_b_19_66024 = net_66024;
  assign seg_16_16_sp4_v_b_2_62066 = net_62066;
  assign seg_16_16_sp4_v_b_34_62320 = net_62320;
  assign seg_16_16_sp4_v_t_36_62555 = seg_15_20_sp4_r_v_b_1_62555;
  assign seg_16_16_sp4_v_t_47_62566 = seg_15_19_sp4_r_v_b_23_62566;
  assign seg_16_17_lutff_1_out_62409 = net_62409;
  assign seg_16_17_sp4_h_l_40_51059 = seg_13_17_sp4_h_r_16_51059;
  assign seg_16_17_sp4_h_l_44_51063 = seg_13_17_sp4_h_r_20_51063;
  assign seg_16_17_sp4_h_l_46_51055 = seg_13_17_sp4_h_r_22_51055;
  assign seg_16_17_sp4_h_l_47_51054 = seg_12_17_sp4_h_r_10_51054;
  assign seg_16_17_sp4_v_b_2_62189 = seg_16_15_sp4_v_b_26_62189;
  assign seg_16_18_lutff_2_out_62533 = net_62533;
  assign seg_16_18_lutff_3_out_62534 = net_62534;
  assign seg_16_18_lutff_4_out_62535 = net_62535;
  assign seg_16_18_neigh_op_lft_2_58703 = seg_15_18_lutff_2_out_58703;
  assign seg_16_18_neigh_op_tnl_3_58827 = seg_15_19_lutff_3_out_58827;
  assign seg_16_18_neigh_op_top_5_62659 = seg_16_19_lutff_5_out_62659;
  assign seg_16_18_sp4_h_l_37_51175 = seg_12_18_sp4_h_r_0_51175;
  assign seg_16_18_sp4_h_r_1_66498 = seg_17_18_sp4_h_r_12_66498;
  assign seg_16_18_sp4_h_r_4_66503 = net_66503;
  assign seg_16_18_sp4_v_t_37_62802 = seg_15_21_sp4_r_v_b_13_62802;
  assign seg_16_19_lutff_1_out_62655 = net_62655;
  assign seg_16_19_lutff_3_out_62657 = net_62657;
  assign seg_16_19_lutff_4_out_62658 = net_62658;
  assign seg_16_19_lutff_5_out_62659 = net_62659;
  assign seg_16_19_lutff_6_out_62660 = net_62660;
  assign seg_16_19_lutff_7_out_62661 = net_62661;
  assign seg_16_19_neigh_op_top_2_62779 = seg_16_20_lutff_2_out_62779;
  assign seg_16_19_neigh_op_top_7_62784 = seg_16_20_lutff_7_out_62784;
  assign seg_16_19_sp4_h_l_41_51304 = seg_12_19_sp4_h_r_4_51304;
  assign seg_16_19_sp4_h_l_42_51307 = seg_13_19_sp4_h_r_18_51307;
  assign seg_16_20_lutff_1_out_62778 = net_62778;
  assign seg_16_20_lutff_2_out_62779 = net_62779;
  assign seg_16_20_lutff_3_out_62780 = net_62780;
  assign seg_16_20_lutff_4_out_62781 = net_62781;
  assign seg_16_20_lutff_5_out_62782 = net_62782;
  assign seg_16_20_lutff_7_out_62784 = net_62784;
  assign seg_16_20_neigh_op_rgt_2_66610 = seg_17_20_lutff_2_out_66610;
  assign seg_16_20_neigh_op_top_7_62907 = seg_16_21_lutff_7_out_62907;
  assign seg_16_20_sp4_h_l_44_51432 = seg_15_20_sp4_h_r_44_51432;
  assign seg_16_20_sp4_v_b_10_62566 = seg_15_19_sp4_r_v_b_23_62566;
  assign seg_16_21_lutff_7_out_62907 = net_62907;
  assign seg_16_21_sp4_h_l_37_51544 = seg_12_21_sp4_h_r_0_51544;
  assign seg_16_21_sp4_h_l_41_51550 = seg_12_21_sp4_h_r_4_51550;
  assign seg_16_21_sp4_h_l_44_51555 = seg_15_21_sp4_h_r_44_51555;
  assign seg_16_21_sp4_v_t_46_63180 = seg_15_25_sp4_r_v_b_11_63180;
  assign seg_16_23_sp4_h_l_42_51799 = seg_15_23_sp4_h_r_42_51799;
  assign seg_16_23_sp4_v_t_38_63418 = seg_15_25_sp4_r_v_b_27_63418;
  assign seg_16_28_lutff_1_out_63762 = net_63762;
  assign seg_16_28_lutff_2_out_63763 = net_63763;
  assign seg_16_28_lutff_3_out_63764 = net_63764;
  assign seg_16_28_lutff_5_out_63766 = net_63766;
  assign seg_16_28_lutff_6_out_63767 = net_63767;
  assign seg_16_28_lutff_7_out_63768 = net_63768;
  assign seg_16_28_neigh_op_top_0_63884 = seg_16_29_lutff_0_out_63884;
  assign seg_16_28_neigh_op_top_4_63888 = seg_16_29_lutff_4_out_63888;
  assign seg_16_28_sp4_v_b_8_63548 = net_63548;
  assign seg_16_29_lutff_0_out_63884 = net_63884;
  assign seg_16_29_lutff_2_out_63886 = net_63886;
  assign seg_16_29_lutff_4_out_63888 = net_63888;
  assign seg_16_29_lutff_6_out_63890 = net_63890;
  assign seg_16_29_neigh_op_bot_1_63762 = seg_16_28_lutff_1_out_63762;
  assign seg_16_29_neigh_op_bot_3_63764 = seg_16_28_lutff_3_out_63764;
  assign seg_16_29_neigh_op_bot_5_63766 = seg_16_28_lutff_5_out_63766;
  assign seg_16_29_neigh_op_bot_6_63767 = seg_16_28_lutff_6_out_63767;
  assign seg_16_29_sp4_r_v_b_32_67748 = seg_17_31_span4_vert_8_67748;
  assign seg_16_2_lutff_1_out_60528 = net_60528;
  assign seg_16_2_lutff_2_out_60529 = net_60529;
  assign seg_16_2_lutff_5_out_60532 = net_60532;
  assign seg_16_2_neigh_op_lft_0_56697 = seg_15_2_lutff_0_out_56697;
  assign seg_16_2_neigh_op_lft_1_56698 = seg_15_2_lutff_1_out_56698;
  assign seg_16_2_neigh_op_lft_6_56703 = seg_15_2_lutff_6_out_56703;
  assign seg_16_2_neigh_op_tnl_7_56863 = seg_15_3_lutff_7_out_56863;
  assign seg_16_31_span4_vert_7_63914 = seg_15_29_sp4_r_v_b_31_63914;
  assign seg_16_5_lutff_2_out_60934 = net_60934;
  assign seg_16_5_lutff_3_out_60935 = net_60935;
  assign seg_16_5_lutff_4_out_60936 = net_60936;
  assign seg_16_5_lutff_5_out_60937 = net_60937;
  assign seg_16_5_lutff_6_out_60938 = net_60938;
  assign seg_16_5_lutff_7_out_60939 = net_60939;
  assign seg_16_5_neigh_op_rgt_0_64763 = seg_17_5_lutff_0_out_64763;
  assign seg_16_5_neigh_op_rgt_1_64764 = seg_17_5_lutff_1_out_64764;
  assign seg_16_5_neigh_op_rgt_2_64765 = seg_17_5_lutff_2_out_64765;
  assign seg_16_5_neigh_op_rgt_3_64766 = seg_17_5_lutff_3_out_64766;
  assign seg_16_5_neigh_op_rgt_6_64769 = seg_17_5_lutff_6_out_64769;
  assign seg_16_5_neigh_op_rgt_7_64770 = seg_17_5_lutff_7_out_64770;
  assign seg_16_5_sp4_h_r_18_61076 = seg_18_5_sp4_h_r_42_61076;
  assign seg_16_6_lutff_0_out_61055 = net_61055;
  assign seg_16_6_neigh_op_rgt_0_64886 = seg_17_6_lutff_0_out_64886;
  assign seg_16_6_sp4_h_l_36_49700 = seg_15_6_sp4_h_r_36_49700;
  assign seg_16_6_sp4_h_r_6_65029 = seg_18_6_sp4_h_r_30_65029;
  assign seg_16_6_sp4_v_b_6_60840 = seg_15_3_sp4_r_v_b_43_60840;
  assign seg_16_7_sp4_v_b_8_60965 = seg_15_6_sp4_r_v_b_21_60965;
  assign seg_16_9_lutff_2_out_61426 = net_61426;
  assign seg_16_9_lutff_3_out_61427 = net_61427;
  assign seg_16_9_lutff_4_out_61428 = net_61428;
  assign seg_16_9_lutff_5_out_61429 = net_61429;
  assign seg_16_9_lutff_6_out_61430 = net_61430;
  assign seg_16_9_sp12_v_b_14_64773 = net_64773;
  assign seg_16_9_sp4_v_b_0_61203 = seg_15_6_sp4_r_v_b_37_61203;
  assign seg_16_9_sp4_v_b_36_61571 = net_61571;
  assign seg_16_9_sp4_v_b_44_61579 = net_61579;
  assign seg_16_9_sp4_v_b_4_61207 = seg_15_8_sp4_r_v_b_17_61207;
  assign seg_17_0_span12_vert_16_68077 = net_68077;
  assign seg_17_0_span4_horz_r_0_68093 = seg_18_0_span4_horz_r_4_68093;
  assign seg_17_0_span4_vert_16_64390 = net_64390;
  assign seg_17_0_span4_vert_18_64392 = net_64392;
  assign seg_17_10_sp4_h_l_37_54022 = seg_15_10_sp4_h_r_24_54022;
  assign seg_17_10_sp4_h_r_11_69347 = seg_18_10_sp4_h_r_22_69347;
  assign seg_17_11_sp4_v_b_10_65290 = seg_17_9_sp4_v_b_34_65290;
  assign seg_17_12_sp4_h_l_37_54268 = seg_13_12_sp4_h_r_0_54268;
  assign seg_17_12_sp4_h_r_18_65768 = net_65768;
  assign seg_17_12_sp4_v_t_39_65897 = seg_16_15_sp4_r_v_b_15_65897;
  assign seg_17_13_lutff_3_out_65750 = net_65750;
  assign seg_17_13_neigh_op_lft_0_61916 = seg_16_13_lutff_0_out_61916;
  assign seg_17_13_neigh_op_lft_3_61919 = seg_16_13_lutff_3_out_61919;
  assign seg_17_13_sp4_h_r_0_69713 = seg_19_13_sp4_h_r_24_69713;
  assign seg_17_13_sp4_h_r_20_65893 = seg_19_13_sp4_h_r_44_65893;
  assign seg_17_13_sp4_r_v_b_29_69606 = net_69606;
  assign seg_17_13_sp4_v_t_43_66024 = seg_16_16_sp4_r_v_b_19_66024;
  assign seg_17_14_lutff_0_out_65870 = net_65870;
  assign seg_17_14_lutff_2_out_65872 = net_65872;
  assign seg_17_14_lutff_3_out_65873 = net_65873;
  assign seg_17_14_lutff_4_out_65874 = net_65874;
  assign seg_17_14_lutff_5_out_65875 = net_65875;
  assign seg_17_14_lutff_7_out_65877 = net_65877;
  assign seg_17_14_neigh_op_top_0_65993 = seg_17_15_lutff_0_out_65993;
  assign seg_17_14_sp4_h_l_37_54514 = seg_13_14_sp4_h_r_0_54514;
  assign seg_17_14_sp4_h_l_38_54519 = seg_14_14_sp4_h_r_14_54519;
  assign seg_17_14_sp4_h_l_44_54525 = seg_14_14_sp4_h_r_20_54525;
  assign seg_17_14_sp4_h_r_26_62178 = seg_15_14_sp4_h_r_2_62178;
  assign seg_17_14_sp4_r_v_b_27_69727 = net_69727;
  assign seg_17_14_sp4_v_b_11_65658 = seg_16_12_sp4_r_v_b_35_65658;
  assign seg_17_15_lutff_0_out_65993 = net_65993;
  assign seg_17_15_lutff_4_out_65997 = net_65997;
  assign seg_17_15_neigh_op_bot_0_65870 = seg_17_14_lutff_0_out_65870;
  assign seg_17_15_sp4_h_l_37_54637 = seg_13_15_sp4_h_r_0_54637;
  assign seg_17_15_sp4_h_r_16_66135 = seg_19_15_sp4_h_r_40_66135;
  assign seg_17_15_sp4_h_r_6_69967 = net_69967;
  assign seg_17_15_sp4_r_v_b_5_69606 = seg_17_13_sp4_r_v_b_29_69606;
  assign seg_17_16_lutff_1_out_66117 = net_66117;
  assign seg_17_16_sp4_h_r_14_66256 = net_66256;
  assign seg_17_16_sp4_h_r_30_62428 = net_62428;
  assign seg_17_16_sp4_v_b_8_65903 = seg_16_15_sp4_r_v_b_21_65903;
  assign seg_17_17_lutff_0_out_66239 = net_66239;
  assign seg_17_17_lutff_2_out_66241 = net_66241;
  assign seg_17_17_neigh_op_bnl_1_62286 = seg_16_16_lutff_1_out_62286;
  assign seg_17_17_neigh_op_bot_1_66117 = seg_17_16_lutff_1_out_66117;
  assign seg_17_17_neigh_op_lft_1_62409 = seg_16_17_lutff_1_out_62409;
  assign seg_17_17_neigh_op_top_2_66364 = seg_17_18_lutff_2_out_66364;
  assign seg_17_17_sp4_h_r_10_70207 = net_70207;
  assign seg_17_17_sp4_h_r_14_66379 = net_66379;
  assign seg_17_17_sp4_h_r_2_70209 = net_70209;
  assign seg_17_17_sp4_v_t_42_66515 = seg_17_20_sp4_v_b_18_66515;
  assign seg_17_18_lutff_0_out_66362 = net_66362;
  assign seg_17_18_lutff_1_out_66363 = net_66363;
  assign seg_17_18_lutff_2_out_66364 = net_66364;
  assign seg_17_18_lutff_4_out_66366 = net_66366;
  assign seg_17_18_neigh_op_lft_2_62533 = seg_16_18_lutff_2_out_62533;
  assign seg_17_18_neigh_op_top_6_66491 = seg_17_19_lutff_6_out_66491;
  assign seg_17_18_sp12_h_r_4_62662 = net_62662;
  assign seg_17_18_sp4_h_l_38_55011 = seg_14_18_sp4_h_r_14_55011;
  assign seg_17_18_sp4_h_r_12_66498 = net_66498;
  assign seg_17_18_sp4_h_r_14_66502 = net_66502;
  assign seg_17_18_sp4_h_r_22_66500 = net_66500;
  assign seg_17_18_sp4_h_r_36_58837 = seg_15_18_sp4_h_r_12_58837;
  assign seg_17_18_sp4_h_r_44_58847 = net_58847;
  assign seg_17_18_sp4_r_v_b_45_70349 = net_70349;
  assign seg_17_18_sp4_v_b_44_66517 = net_66517;
  assign seg_17_19_lutff_1_out_66486 = net_66486;
  assign seg_17_19_lutff_5_out_66490 = net_66490;
  assign seg_17_19_lutff_6_out_66491 = net_66491;
  assign seg_17_19_lutff_7_out_66492 = net_66492;
  assign seg_17_19_neigh_op_lft_1_62655 = seg_16_19_lutff_1_out_62655;
  assign seg_17_19_neigh_op_lft_6_62660 = seg_16_19_lutff_6_out_62660;
  assign seg_17_19_neigh_op_tnl_3_62780 = seg_16_20_lutff_3_out_62780;
  assign seg_17_19_neigh_op_top_0_66608 = seg_17_20_lutff_0_out_66608;
  assign seg_17_19_sp4_h_l_39_55133 = seg_13_19_sp4_h_r_2_55133;
  assign seg_17_19_sp4_h_l_45_55139 = seg_13_19_sp4_h_r_8_55139;
  assign seg_17_19_sp4_h_r_24_62789 = net_62789;
  assign seg_17_19_sp4_h_r_30_62797 = seg_15_19_sp4_h_r_6_62797;
  assign seg_17_19_sp4_h_r_8_70461 = net_70461;
  assign seg_17_19_sp4_r_v_b_29_70344 = net_70344;
  assign seg_17_20_lutff_0_out_66608 = net_66608;
  assign seg_17_20_lutff_1_out_66609 = net_66609;
  assign seg_17_20_lutff_2_out_66610 = net_66610;
  assign seg_17_20_lutff_5_out_66613 = net_66613;
  assign seg_17_20_lutff_6_out_66614 = net_66614;
  assign seg_17_20_neigh_op_lft_5_62782 = seg_16_20_lutff_5_out_62782;
  assign seg_17_20_neigh_op_top_6_66737 = seg_17_21_lutff_6_out_66737;
  assign seg_17_20_sp4_v_b_18_66515 = net_66515;
  assign seg_17_21_lutff_6_out_66737 = net_66737;
  assign seg_17_21_sp4_h_l_41_55381 = seg_15_21_sp4_h_r_28_55381;
  assign seg_17_21_sp4_r_v_b_11_70350 = net_70350;
  assign seg_17_21_sp4_v_b_9_66517 = seg_17_18_sp4_v_b_44_66517;
  assign seg_17_29_neigh_op_bnl_1_63762 = seg_16_28_lutff_1_out_63762;
  assign seg_17_29_neigh_op_bnl_3_63764 = seg_16_28_lutff_3_out_63764;
  assign seg_17_29_neigh_op_bnl_5_63766 = seg_16_28_lutff_5_out_63766;
  assign seg_17_29_neigh_op_bnl_6_63767 = seg_16_28_lutff_6_out_63767;
  assign seg_17_29_sp4_r_v_b_29_71574 = net_71574;
  assign seg_17_2_sp4_v_b_5_64390 = seg_17_0_span4_vert_16_64390;
  assign seg_17_2_sp4_v_b_7_64392 = seg_17_0_span4_vert_18_64392;
  assign seg_17_31_span4_vert_8_67748 = net_67748;
  assign seg_17_5_lutff_0_out_64763 = net_64763;
  assign seg_17_5_lutff_1_out_64764 = net_64764;
  assign seg_17_5_lutff_2_out_64765 = net_64765;
  assign seg_17_5_lutff_3_out_64766 = net_64766;
  assign seg_17_5_lutff_5_out_64768 = net_64768;
  assign seg_17_5_lutff_6_out_64769 = net_64769;
  assign seg_17_5_lutff_7_out_64770 = net_64770;
  assign seg_17_5_neigh_op_lft_2_60934 = seg_16_5_lutff_2_out_60934;
  assign seg_17_5_neigh_op_lft_3_60935 = seg_16_5_lutff_3_out_60935;
  assign seg_17_5_neigh_op_lft_4_60936 = seg_16_5_lutff_4_out_60936;
  assign seg_17_5_neigh_op_lft_5_60937 = seg_16_5_lutff_5_out_60937;
  assign seg_17_5_neigh_op_lft_6_60938 = seg_16_5_lutff_6_out_60938;
  assign seg_17_5_neigh_op_lft_7_60939 = seg_16_5_lutff_7_out_60939;
  assign seg_17_5_neigh_op_tnr_0_68717 = seg_18_6_lutff_0_out_68717;
  assign seg_17_6_lutff_0_out_64886 = net_64886;
  assign seg_17_6_lutff_4_out_64890 = net_64890;
  assign seg_17_6_lutff_5_out_64891 = net_64891;
  assign seg_17_6_lutff_7_out_64893 = net_64893;
  assign seg_17_6_neigh_op_bnr_5_68599 = seg_18_5_lutff_5_out_68599;
  assign seg_17_6_neigh_op_bot_1_64764 = seg_17_5_lutff_1_out_64764;
  assign seg_17_6_neigh_op_bot_2_64765 = seg_17_5_lutff_2_out_64765;
  assign seg_17_6_neigh_op_bot_6_64769 = seg_17_5_lutff_6_out_64769;
  assign seg_17_6_neigh_op_bot_7_64770 = seg_17_5_lutff_7_out_64770;
  assign seg_17_6_neigh_op_lft_0_61055 = seg_16_6_lutff_0_out_61055;
  assign seg_17_6_neigh_op_rgt_0_68717 = seg_18_6_lutff_0_out_68717;
  assign seg_17_6_neigh_op_rgt_7_68724 = seg_18_6_lutff_7_out_68724;
  assign seg_17_9_lutff_1_out_65256 = net_65256;
  assign seg_17_9_sp12_v_b_0_68077 = seg_17_0_span12_vert_16_68077;
  assign seg_17_9_sp4_v_b_34_65290 = net_65290;
  assign seg_18_0_span4_horz_r_4_68093 = net_68093;
  assign seg_18_10_sp4_h_l_44_57863 = seg_15_10_sp4_h_r_20_57863;
  assign seg_18_10_sp4_h_r_22_69347 = net_69347;
  assign seg_18_10_sp4_h_r_38_61687 = net_61687;
  assign seg_18_10_sp4_h_r_6_73183 = net_73183;
  assign seg_18_10_sp4_v_b_22_69120 = net_69120;
  assign seg_18_11_sp4_h_l_41_57981 = seg_14_11_sp4_h_r_4_57981;
  assign seg_18_12_sp4_h_r_12_69591 = net_69591;
  assign seg_18_12_sp4_h_r_30_65767 = net_65767;
  assign seg_18_12_sp4_h_r_6_73429 = net_73429;
  assign seg_18_13_lutff_1_out_69579 = net_69579;
  assign seg_18_13_neigh_op_lft_3_65750 = seg_17_13_lutff_3_out_65750;
  assign seg_18_13_neigh_op_top_4_69705 = seg_18_14_lutff_4_out_69705;
  assign seg_18_13_sp12_h_r_4_65878 = net_65878;
  assign seg_18_13_sp4_h_l_36_58222 = seg_15_13_sp4_h_r_12_58222;
  assign seg_18_13_sp4_h_l_39_58225 = seg_14_13_sp4_h_r_2_58225;
  assign seg_18_13_sp4_h_l_42_58230 = seg_15_13_sp4_h_r_18_58230;
  assign seg_18_13_sp4_h_l_43_58229 = seg_14_13_sp4_h_r_6_58229;
  assign seg_18_13_sp4_h_l_45_58231 = seg_14_13_sp4_h_r_8_58231;
  assign seg_18_13_sp4_h_l_47_58223 = seg_14_13_sp4_h_r_10_58223;
  assign seg_18_13_sp4_h_r_0_73544 = net_73544;
  assign seg_18_13_sp4_h_r_10_73546 = seg_20_13_sp4_h_r_34_73546;
  assign seg_18_13_sp4_h_r_12_69714 = seg_20_13_sp4_h_r_36_69714;
  assign seg_18_13_sp4_h_r_14_69718 = net_69718;
  assign seg_18_13_sp4_h_r_22_69716 = net_69716;
  assign seg_18_13_sp4_h_r_26_65886 = net_65886;
  assign seg_18_13_sp4_h_r_41_62057 = seg_15_13_sp4_h_r_4_62057;
  assign seg_18_13_sp4_h_r_47_62053 = seg_15_13_sp4_h_r_10_62053;
  assign seg_18_13_sp4_h_r_4_73550 = net_73550;
  assign seg_18_13_sp4_h_r_8_73554 = net_73554;
  assign seg_18_14_lutff_1_out_69702 = net_69702;
  assign seg_18_14_lutff_4_out_69705 = net_69705;
  assign seg_18_14_lutff_7_out_69708 = net_69708;
  assign seg_18_14_neigh_op_bnr_1_73410 = seg_19_13_ram_RDATA_14_73410;
  assign seg_18_14_neigh_op_bnr_7_73416 = seg_19_13_ram_RDATA_8_73416;
  assign seg_18_14_neigh_op_bot_1_69579 = seg_18_13_lutff_1_out_69579;
  assign seg_18_14_neigh_op_lft_2_65872 = seg_17_14_lutff_2_out_65872;
  assign seg_18_14_neigh_op_lft_3_65873 = seg_17_14_lutff_3_out_65873;
  assign seg_18_14_neigh_op_lft_4_65874 = seg_17_14_lutff_4_out_65874;
  assign seg_18_14_neigh_op_lft_7_65877 = seg_17_14_lutff_7_out_65877;
  assign seg_18_14_neigh_op_tnr_2_73657 = seg_19_15_ram_RDATA_13_73657;
  assign seg_18_14_neigh_op_tnr_5_73660 = seg_19_15_ram_RDATA_10_73660;
  assign seg_18_14_sp4_h_l_37_58344 = seg_14_14_sp4_h_r_0_58344;
  assign seg_18_14_sp4_h_l_38_58349 = seg_15_14_sp4_h_r_14_58349;
  assign seg_18_14_sp4_h_r_0_73667 = net_73667;
  assign seg_18_14_sp4_h_r_10_73669 = net_73669;
  assign seg_18_14_sp4_h_r_20_69847 = net_69847;
  assign seg_18_14_sp4_h_r_6_73675 = net_73675;
  assign seg_18_14_sp4_r_v_b_38_73681 = seg_19_16_sp4_v_b_14_73681;
  assign seg_18_15_sp4_h_r_0_73790 = net_73790;
  assign seg_18_15_sp4_h_r_14_69964 = net_69964;
  assign seg_18_15_sp4_h_r_20_69970 = net_69970;
  assign seg_18_15_sp4_h_r_28_66134 = seg_16_15_sp4_h_r_4_66134;
  assign seg_18_15_sp4_h_r_34_66130 = seg_16_15_sp4_h_r_10_66130;
  assign seg_18_15_sp4_h_r_40_62304 = net_62304;
  assign seg_18_15_sp4_h_r_41_62303 = seg_15_15_sp4_h_r_4_62303;
  assign seg_18_15_sp4_h_r_44_62308 = net_62308;
  assign seg_18_15_sp4_h_r_45_62307 = seg_15_15_sp4_h_r_8_62307;
  assign seg_18_15_sp4_r_v_b_11_73443 = net_73443;
  assign seg_18_15_sp4_r_v_b_7_73439 = net_73439;
  assign seg_18_16_lutff_2_out_69949 = net_69949;
  assign seg_18_16_sp4_h_r_20_70093 = net_70093;
  assign seg_18_16_sp4_h_r_4_73919 = net_73919;
  assign seg_18_16_sp4_r_v_b_37_73926 = net_73926;
  assign seg_18_16_sp4_r_v_b_5_73560 = net_73560;
  assign seg_18_16_sp4_v_b_3_69727 = seg_17_14_sp4_r_v_b_27_69727;
  assign seg_18_17_neigh_op_lft_0_66239 = seg_17_17_lutff_0_out_66239;
  assign seg_18_17_neigh_op_top_4_70197 = seg_18_18_lutff_4_out_70197;
  assign seg_18_17_sp4_h_r_0_74036 = net_74036;
  assign seg_18_17_sp4_h_r_10_74038 = net_74038;
  assign seg_18_17_sp4_h_r_12_70206 = net_70206;
  assign seg_18_17_sp4_h_r_2_74040 = net_74040;
  assign seg_18_17_sp4_h_r_30_66382 = net_66382;
  assign seg_18_17_sp4_h_r_38_62548 = net_62548;
  assign seg_18_17_sp4_h_r_4_74042 = net_74042;
  assign seg_18_17_sp4_h_r_8_74046 = net_74046;
  assign seg_18_17_sp4_h_r_9_74047 = seg_21_17_sp4_h_r_44_74047;
  assign seg_18_17_sp4_v_t_40_70344 = seg_17_19_sp4_r_v_b_29_70344;
  assign seg_18_17_sp4_v_t_46_70350 = seg_17_21_sp4_r_v_b_11_70350;
  assign seg_18_18_lutff_3_out_70196 = net_70196;
  assign seg_18_18_lutff_4_out_70197 = net_70197;
  assign seg_18_18_lutff_5_out_70198 = net_70198;
  assign seg_18_18_neigh_op_bnr_7_73908 = seg_19_17_ram_RDATA_8_73908;
  assign seg_18_18_neigh_op_lft_0_66362 = seg_17_18_lutff_0_out_66362;
  assign seg_18_18_neigh_op_lft_1_66363 = seg_17_18_lutff_1_out_66363;
  assign seg_18_18_neigh_op_lft_4_66366 = seg_17_18_lutff_4_out_66366;
  assign seg_18_18_neigh_op_rgt_1_74025 = seg_19_18_ram_RDATA_6_74025;
  assign seg_18_18_neigh_op_rgt_2_74026 = seg_19_18_ram_RDATA_5_74026;
  assign seg_18_18_neigh_op_rgt_5_74029 = seg_19_18_ram_RDATA_2_74029;
  assign seg_18_18_neigh_op_top_7_70323 = seg_18_19_lutff_7_out_70323;
  assign seg_18_18_sp12_h_r_3_70324 = seg_21_18_sp12_h_r_8_70324;
  assign seg_18_18_sp4_h_l_36_58837 = seg_15_18_sp4_h_r_12_58837;
  assign seg_18_18_sp4_h_l_45_58846 = seg_14_18_sp4_h_r_8_58846;
  assign seg_18_18_sp4_h_r_12_70329 = net_70329;
  assign seg_18_18_sp4_h_r_27_66502 = seg_17_18_sp4_h_r_14_66502;
  assign seg_18_18_sp4_h_r_30_66505 = net_66505;
  assign seg_18_18_sp4_h_r_4_74165 = net_74165;
  assign seg_18_19_lutff_7_out_70323 = net_70323;
  assign seg_18_19_sp4_h_l_46_58962 = seg_15_19_sp4_h_r_22_58962;
  assign seg_18_20_neigh_op_lft_1_66609 = seg_17_20_lutff_1_out_66609;
  assign seg_18_20_sp4_h_l_47_59084 = seg_14_20_sp4_h_r_10_59084;
  assign seg_18_20_sp4_r_v_b_31_74300 = net_74300;
  assign seg_18_21_sp4_v_b_8_70349 = seg_17_18_sp4_r_v_b_45_70349;
  assign seg_18_27_sp4_v_t_41_71575 = seg_18_31_span4_vert_4_71575;
  assign seg_18_27_sp4_v_t_43_71577 = seg_18_31_span4_vert_6_71577;
  assign seg_18_2_sp4_h_l_47_56870 = seg_14_2_sp4_h_r_10_56870;
  assign seg_18_30_sp4_v_t_36_75655 = seg_18_31_span4_vert_36_75655;
  assign seg_18_31_span4_vert_36_75655 = net_75655;
  assign seg_18_31_span4_vert_4_71575 = net_71575;
  assign seg_18_31_span4_vert_5_71574 = seg_17_29_sp4_r_v_b_29_71574;
  assign seg_18_31_span4_vert_6_71577 = net_71577;
  assign seg_18_5_lutff_5_out_68599 = net_68599;
  assign seg_18_5_lutff_7_out_68601 = net_68601;
  assign seg_18_5_neigh_op_top_0_68717 = seg_18_6_lutff_0_out_68717;
  assign seg_18_5_sp4_h_r_42_61076 = net_61076;
  assign seg_18_6_lutff_0_out_68717 = net_68717;
  assign seg_18_6_lutff_2_out_68719 = net_68719;
  assign seg_18_6_lutff_5_out_68722 = net_68722;
  assign seg_18_6_lutff_7_out_68724 = net_68724;
  assign seg_18_6_neigh_op_bnl_5_64768 = seg_17_5_lutff_5_out_64768;
  assign seg_18_6_neigh_op_bot_5_68599 = seg_18_5_lutff_5_out_68599;
  assign seg_18_6_neigh_op_lft_4_64890 = seg_17_6_lutff_4_out_64890;
  assign seg_18_6_neigh_op_lft_5_64891 = seg_17_6_lutff_5_out_64891;
  assign seg_18_6_neigh_op_lft_7_64893 = seg_17_6_lutff_7_out_64893;
  assign seg_18_6_sp4_h_r_10_72685 = net_72685;
  assign seg_18_6_sp4_h_r_2_72687 = net_72687;
  assign seg_18_6_sp4_h_r_30_65029 = net_65029;
  assign seg_18_6_sp4_h_r_44_61201 = net_61201;
  assign seg_18_6_sp4_h_r_7_72692 = seg_21_6_sp4_h_r_42_72692;
  assign seg_18_7_sp4_v_t_46_69120 = seg_18_10_sp4_v_b_22_69120;
  assign seg_18_8_sp4_h_l_45_57616 = seg_14_8_sp4_h_r_8_57616;
  assign seg_19_10_sp4_h_r_0_76795 = seg_21_10_sp4_h_r_24_76795;
  assign seg_19_10_sp4_h_r_10_76797 = seg_21_10_sp4_h_r_34_76797;
  assign seg_19_10_sp4_h_r_3_76800 = seg_20_10_sp4_h_r_14_76800;
  assign seg_19_12_sp4_h_l_36_61929 = seg_16_12_sp4_h_r_12_61929;
  assign seg_19_12_sp4_v_t_43_73563 = seg_19_16_sp4_v_b_6_73563;
  assign seg_19_13_ram_RDATA_10_73414 = net_73414;
  assign seg_19_13_ram_RDATA_12_73412 = net_73412;
  assign seg_19_13_ram_RDATA_13_73411 = net_73411;
  assign seg_19_13_ram_RDATA_14_73410 = net_73410;
  assign seg_19_13_ram_RDATA_8_73416 = net_73416;
  assign seg_19_13_sp4_h_l_37_62051 = seg_15_13_sp4_h_r_0_62051;
  assign seg_19_13_sp4_h_l_41_62057 = seg_15_13_sp4_h_r_4_62057;
  assign seg_19_13_sp4_h_l_47_62053 = seg_15_13_sp4_h_r_10_62053;
  assign seg_19_13_sp4_h_r_0_77101 = net_77101;
  assign seg_19_13_sp4_h_r_24_69713 = net_69713;
  assign seg_19_13_sp4_h_r_41_65888 = seg_16_13_sp4_h_r_4_65888;
  assign seg_19_13_sp4_h_r_44_65893 = net_65893;
  assign seg_19_14_ram_RDATA_1_73538 = net_73538;
  assign seg_19_14_ram_RDATA_2_73537 = net_73537;
  assign seg_19_14_ram_RDATA_5_73534 = net_73534;
  assign seg_19_14_sp4_h_l_45_62184 = seg_15_14_sp4_h_r_8_62184;
  assign seg_19_14_sp4_h_r_16_73674 = net_73674;
  assign seg_19_14_sp4_h_r_3_77208 = seg_22_14_sp4_h_r_38_77208;
  assign seg_19_14_sp4_r_v_b_26_77116 = seg_20_16_sp4_v_b_2_77116;
  assign seg_19_14_sp4_r_v_b_30_77120 = seg_20_16_sp4_v_b_6_77120;
  assign seg_19_14_sp4_r_v_b_32_77122 = seg_20_16_sp4_v_b_8_77122;
  assign seg_19_14_sp4_r_v_b_34_77124 = seg_20_16_sp4_v_b_10_77124;
  assign seg_19_14_sp4_r_v_b_38_77217 = seg_20_16_sp4_v_b_14_77217;
  assign seg_19_14_sp4_r_v_b_3_76911 = net_76911;
  assign seg_19_14_sp4_r_v_b_41_77220 = net_77220;
  assign seg_19_14_sp4_r_v_b_44_77223 = seg_20_16_sp4_v_b_20_77223;
  assign seg_19_14_sp4_r_v_b_47_77226 = net_77226;
  assign seg_19_14_sp4_r_v_b_7_76915 = net_76915;
  assign seg_19_14_sp4_v_b_29_73560 = seg_18_16_sp4_r_v_b_5_73560;
  assign seg_19_15_ram_RDATA_10_73660 = net_73660;
  assign seg_19_15_ram_RDATA_12_73658 = net_73658;
  assign seg_19_15_ram_RDATA_13_73657 = net_73657;
  assign seg_19_15_ram_RDATA_14_73656 = net_73656;
  assign seg_19_15_ram_RDATA_15_73655 = net_73655;
  assign seg_19_15_sp4_h_l_36_62298 = seg_16_15_sp4_h_r_12_62298;
  assign seg_19_15_sp4_h_l_40_62304 = seg_18_15_sp4_h_r_40_62304;
  assign seg_19_15_sp4_h_l_41_62303 = seg_15_15_sp4_h_r_4_62303;
  assign seg_19_15_sp4_h_l_44_62308 = seg_18_15_sp4_h_r_44_62308;
  assign seg_19_15_sp4_h_l_45_62307 = seg_15_15_sp4_h_r_8_62307;
  assign seg_19_15_sp4_h_r_14_73795 = net_73795;
  assign seg_19_15_sp4_h_r_40_66135 = net_66135;
  assign seg_19_15_sp4_r_v_b_13_77114 = net_77114;
  assign seg_19_15_sp4_v_b_11_73443 = seg_18_15_sp4_r_v_b_11_73443;
  assign seg_19_15_sp4_v_b_7_73439 = seg_18_15_sp4_r_v_b_7_73439;
  assign seg_19_16_neigh_op_lft_2_69949 = seg_18_16_lutff_2_out_69949;
  assign seg_19_16_neigh_op_rgt_1_77264 = seg_20_16_lutff_1_out_77264;
  assign seg_19_16_neigh_op_rgt_2_77265 = seg_20_16_lutff_2_out_77265;
  assign seg_19_16_neigh_op_rgt_3_77266 = seg_20_16_lutff_3_out_77266;
  assign seg_19_16_neigh_op_rgt_4_77267 = seg_20_16_lutff_4_out_77267;
  assign seg_19_16_neigh_op_rgt_5_77268 = seg_20_16_lutff_5_out_77268;
  assign seg_19_16_neigh_op_rgt_6_77269 = seg_20_16_lutff_6_out_77269;
  assign seg_19_16_neigh_op_rgt_7_77270 = seg_20_16_lutff_7_out_77270;
  assign seg_19_16_ram_RDATA_1_73784 = net_73784;
  assign seg_19_16_ram_RDATA_3_73782 = net_73782;
  assign seg_19_16_ram_RDATA_5_73780 = net_73780;
  assign seg_19_16_ram_RDATA_7_73778 = net_73778;
  assign seg_19_16_sp4_h_r_0_77407 = seg_21_16_sp4_h_r_24_77407;
  assign seg_19_16_sp4_h_r_26_70086 = net_70086;
  assign seg_19_16_sp4_r_v_b_19_77222 = net_77222;
  assign seg_19_16_sp4_v_b_14_73681 = net_73681;
  assign seg_19_16_sp4_v_b_6_73563 = net_73563;
  assign seg_19_17_ram_RDATA_10_73906 = net_73906;
  assign seg_19_17_ram_RDATA_11_73905 = net_73905;
  assign seg_19_17_ram_RDATA_12_73904 = net_73904;
  assign seg_19_17_ram_RDATA_8_73908 = net_73908;
  assign seg_19_17_sp4_h_l_38_62548 = seg_18_17_sp4_h_r_38_62548;
  assign seg_19_17_sp4_h_r_0_77509 = net_77509;
  assign seg_19_17_sp4_h_r_11_77512 = seg_22_17_sp4_h_r_46_77512;
  assign seg_19_17_sp4_h_r_1_77510 = seg_22_17_sp4_h_r_36_77510;
  assign seg_19_17_sp4_h_r_26_70209 = seg_17_17_sp4_h_r_2_70209;
  assign seg_19_17_sp4_h_r_28_70211 = net_70211;
  assign seg_19_17_sp4_h_r_2_77513 = net_77513;
  assign seg_19_17_sp4_h_r_34_70207 = seg_17_17_sp4_h_r_10_70207;
  assign seg_19_17_sp4_h_r_3_77514 = seg_22_17_sp4_h_r_38_77514;
  assign seg_19_17_sp4_h_r_5_77516 = seg_22_17_sp4_h_r_40_77516;
  assign seg_19_17_sp4_h_r_7_77518 = seg_22_17_sp4_h_r_42_77518;
  assign seg_19_17_sp4_r_v_b_5_77219 = net_77219;
  assign seg_19_17_sp4_v_t_40_74175 = seg_19_18_sp4_v_b_40_74175;
  assign seg_19_18_ram_RDATA_0_74031 = net_74031;
  assign seg_19_18_ram_RDATA_1_74030 = net_74030;
  assign seg_19_18_ram_RDATA_2_74029 = net_74029;
  assign seg_19_18_ram_RDATA_4_74027 = net_74027;
  assign seg_19_18_ram_RDATA_5_74026 = net_74026;
  assign seg_19_18_ram_RDATA_6_74025 = net_74025;
  assign seg_19_18_ram_RDATA_7_74024 = net_74024;
  assign seg_19_18_sp4_h_l_37_62666 = seg_15_18_sp4_h_r_0_62666;
  assign seg_19_18_sp4_h_r_41_66503 = seg_16_18_sp4_h_r_4_66503;
  assign seg_19_18_sp4_r_v_b_10_77328 = seg_20_16_sp4_v_b_34_77328;
  assign seg_19_18_sp4_r_v_b_14_77421 = seg_20_16_sp4_v_b_38_77421;
  assign seg_19_18_sp4_r_v_b_16_77423 = seg_20_16_sp4_v_b_40_77423;
  assign seg_19_18_sp4_r_v_b_4_77322 = seg_20_16_sp4_v_b_28_77322;
  assign seg_19_18_sp4_v_b_13_73926 = seg_18_16_sp4_r_v_b_37_73926;
  assign seg_19_18_sp4_v_b_40_74175 = net_74175;
  assign seg_19_18_sp4_v_t_42_74300 = seg_18_20_sp4_r_v_b_31_74300;
  assign seg_19_19_sp4_h_l_37_62789 = seg_17_19_sp4_h_r_24_62789;
  assign seg_19_6_sp4_h_l_44_61201 = seg_18_6_sp4_h_r_44_61201;
  assign seg_19_6_sp4_h_r_2_76391 = seg_21_6_sp4_h_r_26_76391;
  assign seg_19_7_sp4_h_r_5_76496 = seg_20_7_sp4_h_r_16_76496;
  assign seg_20_10_lutff_0_out_76651 = net_76651;
  assign seg_20_10_lutff_3_out_76654 = net_76654;
  assign seg_20_10_lutff_7_out_76658 = net_76658;
  assign seg_20_10_neigh_op_bot_1_76550 = seg_20_9_lutff_1_out_76550;
  assign seg_20_10_neigh_op_bot_5_76554 = seg_20_9_lutff_5_out_76554;
  assign seg_20_10_neigh_op_rgt_1_80072 = seg_21_10_lutff_1_out_80072;
  assign seg_20_10_neigh_op_rgt_4_80075 = seg_21_10_lutff_4_out_80075;
  assign seg_20_10_sp12_v_b_14_79589 = net_79589;
  assign seg_20_10_sp4_h_r_0_80206 = net_80206;
  assign seg_20_10_sp4_h_r_10_80208 = net_80208;
  assign seg_20_10_sp4_h_r_14_76800 = net_76800;
  assign seg_20_10_sp4_h_r_7_80215 = seg_21_10_sp4_h_r_18_80215;
  assign seg_20_10_sp4_r_v_b_15_79975 = net_79975;
  assign seg_20_10_sp4_r_v_b_31_80101 = net_80101;
  assign seg_20_10_sp4_r_v_b_47_80229 = net_80229;
  assign seg_20_10_sp4_v_b_46_76817 = net_76817;
  assign seg_20_10_sp4_v_b_6_76508 = net_76508;
  assign seg_20_11_lutff_5_out_76758 = net_76758;
  assign seg_20_12_lutff_0_out_76855 = net_76855;
  assign seg_20_12_lutff_1_out_76856 = net_76856;
  assign seg_20_12_lutff_2_out_76857 = net_76857;
  assign seg_20_12_lutff_3_out_76858 = net_76858;
  assign seg_20_12_lutff_4_out_76859 = net_76859;
  assign seg_20_12_lutff_5_out_76860 = net_76860;
  assign seg_20_12_lutff_6_out_76861 = net_76861;
  assign seg_20_12_lutff_7_out_76862 = net_76862;
  assign seg_20_12_neigh_op_bot_5_76758 = seg_20_11_lutff_5_out_76758;
  assign seg_20_12_neigh_op_rgt_7_80324 = seg_21_12_lutff_7_out_80324;
  assign seg_20_12_neigh_op_tnl_3_73412 = seg_19_13_ram_RDATA_12_73412;
  assign seg_20_12_sp4_h_l_37_65759 = seg_16_12_sp4_h_r_0_65759;
  assign seg_20_12_sp4_h_l_39_65763 = seg_16_12_sp4_h_r_2_65763;
  assign seg_20_12_sp4_h_l_42_65768 = seg_17_12_sp4_h_r_18_65768;
  assign seg_20_12_sp4_h_l_43_65767 = seg_18_12_sp4_h_r_30_65767;
  assign seg_20_12_sp4_h_r_30_73429 = seg_18_12_sp4_h_r_6_73429;
  assign seg_20_12_sp4_h_r_36_69591 = seg_18_12_sp4_h_r_12_69591;
  assign seg_20_12_sp4_r_v_b_10_80106 = seg_21_10_sp4_v_b_34_80106;
  assign seg_20_12_sp4_v_b_27_76911 = seg_19_14_sp4_r_v_b_3_76911;
  assign seg_20_12_sp4_v_b_31_76915 = seg_19_14_sp4_r_v_b_7_76915;
  assign seg_20_12_sp4_v_t_36_77113 = seg_20_15_sp4_v_b_12_77113;
  assign seg_20_13_lutff_0_out_76957 = net_76957;
  assign seg_20_13_lutff_4_out_76961 = net_76961;
  assign seg_20_13_lutff_7_out_76964 = net_76964;
  assign seg_20_13_neigh_op_bot_4_76859 = seg_20_12_lutff_4_out_76859;
  assign seg_20_13_neigh_op_lft_2_73411 = seg_19_13_ram_RDATA_13_73411;
  assign seg_20_13_neigh_op_lft_5_73414 = seg_19_13_ram_RDATA_10_73414;
  assign seg_20_13_neigh_op_tnl_2_73534 = seg_19_14_ram_RDATA_5_73534;
  assign seg_20_13_neigh_op_tnl_5_73537 = seg_19_14_ram_RDATA_2_73537;
  assign seg_20_13_neigh_op_tnl_6_73538 = seg_19_14_ram_RDATA_1_73538;
  assign seg_20_13_neigh_op_top_1_77060 = seg_20_14_lutff_1_out_77060;
  assign seg_20_13_neigh_op_top_2_77061 = seg_20_14_lutff_2_out_77061;
  assign seg_20_13_neigh_op_top_4_77063 = seg_20_14_lutff_4_out_77063;
  assign seg_20_13_neigh_op_top_6_77065 = seg_20_14_lutff_6_out_77065;
  assign seg_20_13_sp12_h_r_8_65878 = seg_18_13_sp12_h_r_4_65878;
  assign seg_20_13_sp4_h_l_39_65886 = seg_18_13_sp4_h_r_26_65886;
  assign seg_20_13_sp4_h_r_28_73550 = seg_18_13_sp4_h_r_4_73550;
  assign seg_20_13_sp4_h_r_34_73546 = net_73546;
  assign seg_20_13_sp4_h_r_36_69714 = net_69714;
  assign seg_20_13_sp4_h_r_38_69718 = seg_18_13_sp4_h_r_14_69718;
  assign seg_20_13_sp4_h_r_42_69722 = net_69722;
  assign seg_20_13_sp4_r_v_b_5_80222 = seg_21_10_sp4_v_b_40_80222;
  assign seg_20_13_sp4_v_b_11_76817 = seg_20_10_sp4_v_b_46_76817;
  assign seg_20_13_sp4_v_b_22_76919 = net_76919;
  assign seg_20_13_sp4_v_b_28_77016 = net_77016;
  assign seg_20_13_sp4_v_b_37_77114 = seg_19_15_sp4_r_v_b_13_77114;
  assign seg_20_13_sp4_v_t_40_77219 = seg_19_17_sp4_r_v_b_5_77219;
  assign seg_20_13_sp4_v_t_41_77220 = seg_19_14_sp4_r_v_b_41_77220;
  assign seg_20_13_sp4_v_t_43_77222 = seg_19_16_sp4_r_v_b_19_77222;
  assign seg_20_13_sp4_v_t_47_77226 = seg_19_14_sp4_r_v_b_47_77226;
  assign seg_20_14_lutff_0_out_77059 = net_77059;
  assign seg_20_14_lutff_1_out_77060 = net_77060;
  assign seg_20_14_lutff_2_out_77061 = net_77061;
  assign seg_20_14_lutff_3_out_77062 = net_77062;
  assign seg_20_14_lutff_4_out_77063 = net_77063;
  assign seg_20_14_lutff_5_out_77064 = net_77064;
  assign seg_20_14_lutff_6_out_77065 = net_77065;
  assign seg_20_14_lutff_7_out_77066 = net_77066;
  assign seg_20_14_neigh_op_bnr_7_80447 = seg_21_13_lutff_7_out_80447;
  assign seg_20_14_neigh_op_bot_7_76964 = seg_20_13_lutff_7_out_76964;
  assign seg_20_14_neigh_op_top_1_77162 = seg_20_15_lutff_1_out_77162;
  assign seg_20_14_sp4_h_r_24_73667 = seg_18_14_sp4_h_r_0_73667;
  assign seg_20_14_sp4_h_r_30_73675 = seg_18_14_sp4_h_r_6_73675;
  assign seg_20_14_sp4_h_r_34_73669 = seg_18_14_sp4_h_r_10_73669;
  assign seg_20_14_sp4_h_r_44_69847 = seg_18_14_sp4_h_r_20_69847;
  assign seg_20_14_sp4_v_b_11_76919 = seg_20_13_sp4_v_b_22_76919;
  assign seg_20_14_sp4_v_b_27_77115 = seg_20_15_sp4_v_b_14_77115;
  assign seg_20_14_sp4_v_t_41_77322 = seg_20_16_sp4_v_b_28_77322;
  assign seg_20_15_lutff_0_out_77161 = net_77161;
  assign seg_20_15_lutff_1_out_77162 = net_77162;
  assign seg_20_15_lutff_2_out_77163 = net_77163;
  assign seg_20_15_lutff_3_out_77164 = net_77164;
  assign seg_20_15_lutff_4_out_77165 = net_77165;
  assign seg_20_15_lutff_5_out_77166 = net_77166;
  assign seg_20_15_neigh_op_lft_0_73655 = seg_19_15_ram_RDATA_15_73655;
  assign seg_20_15_neigh_op_lft_1_73656 = seg_19_15_ram_RDATA_14_73656;
  assign seg_20_15_neigh_op_lft_3_73658 = seg_19_15_ram_RDATA_12_73658;
  assign seg_20_15_neigh_op_tnl_0_73778 = seg_19_16_ram_RDATA_7_73778;
  assign seg_20_15_neigh_op_tnl_2_73780 = seg_19_16_ram_RDATA_5_73780;
  assign seg_20_15_neigh_op_tnl_4_73782 = seg_19_16_ram_RDATA_3_73782;
  assign seg_20_15_neigh_op_tnl_6_73784 = seg_19_16_ram_RDATA_1_73784;
  assign seg_20_15_sp4_h_r_24_73790 = seg_18_15_sp4_h_r_0_73790;
  assign seg_20_15_sp4_h_r_38_69964 = seg_18_15_sp4_h_r_14_69964;
  assign seg_20_15_sp4_h_r_44_69970 = seg_18_15_sp4_h_r_20_69970;
  assign seg_20_15_sp4_v_b_12_77113 = net_77113;
  assign seg_20_15_sp4_v_b_14_77115 = net_77115;
  assign seg_20_15_sp4_v_b_4_77016 = seg_20_13_sp4_v_b_28_77016;
  assign seg_20_16_lutff_1_out_77264 = net_77264;
  assign seg_20_16_lutff_2_out_77265 = net_77265;
  assign seg_20_16_lutff_3_out_77266 = net_77266;
  assign seg_20_16_lutff_4_out_77267 = net_77267;
  assign seg_20_16_lutff_5_out_77268 = net_77268;
  assign seg_20_16_lutff_6_out_77269 = net_77269;
  assign seg_20_16_lutff_7_out_77270 = net_77270;
  assign seg_20_16_sp4_h_r_28_73919 = seg_18_16_sp4_h_r_4_73919;
  assign seg_20_16_sp4_h_r_4_80950 = net_80950;
  assign seg_20_16_sp4_r_v_b_27_80835 = net_80835;
  assign seg_20_16_sp4_r_v_b_31_80839 = net_80839;
  assign seg_20_16_sp4_v_b_10_77124 = net_77124;
  assign seg_20_16_sp4_v_b_14_77217 = net_77217;
  assign seg_20_16_sp4_v_b_20_77223 = net_77223;
  assign seg_20_16_sp4_v_b_28_77322 = net_77322;
  assign seg_20_16_sp4_v_b_2_77116 = net_77116;
  assign seg_20_16_sp4_v_b_34_77328 = net_77328;
  assign seg_20_16_sp4_v_b_38_77421 = net_77421;
  assign seg_20_16_sp4_v_b_40_77423 = net_77423;
  assign seg_20_16_sp4_v_b_6_77120 = net_77120;
  assign seg_20_16_sp4_v_b_8_77122 = net_77122;
  assign seg_20_17_lutff_1_out_77366 = net_77366;
  assign seg_20_17_lutff_2_out_77367 = net_77367;
  assign seg_20_17_lutff_3_out_77368 = net_77368;
  assign seg_20_17_lutff_5_out_77370 = net_77370;
  assign seg_20_17_lutff_6_out_77371 = net_77371;
  assign seg_20_17_lutff_7_out_77372 = net_77372;
  assign seg_20_17_neigh_op_bot_4_77267 = seg_20_16_lutff_4_out_77267;
  assign seg_20_17_neigh_op_bot_5_77268 = seg_20_16_lutff_5_out_77268;
  assign seg_20_17_neigh_op_lft_4_73905 = seg_19_17_ram_RDATA_11_73905;
  assign seg_20_17_neigh_op_rgt_4_80936 = seg_21_17_lutff_4_out_80936;
  assign seg_20_17_neigh_op_rgt_6_80938 = seg_21_17_lutff_6_out_80938;
  assign seg_20_17_neigh_op_tnl_0_74024 = seg_19_18_ram_RDATA_7_74024;
  assign seg_20_17_neigh_op_tnl_6_74030 = seg_19_18_ram_RDATA_1_74030;
  assign seg_20_17_sp12_v_b_1_79589 = seg_20_10_sp12_v_b_14_79589;
  assign seg_20_17_sp4_h_l_38_66379 = seg_17_17_sp4_h_r_14_66379;
  assign seg_20_17_sp4_h_l_43_66382 = seg_18_17_sp4_h_r_30_66382;
  assign seg_20_17_sp4_h_r_1_81068 = seg_21_17_sp4_h_r_12_81068;
  assign seg_20_17_sp4_h_r_26_74040 = seg_18_17_sp4_h_r_2_74040;
  assign seg_20_17_sp4_h_r_32_74046 = seg_18_17_sp4_h_r_8_74046;
  assign seg_20_17_sp4_h_r_36_70206 = seg_18_17_sp4_h_r_12_70206;
  assign seg_20_17_sp4_h_r_41_70211 = seg_19_17_sp4_h_r_28_70211;
  assign seg_20_17_sp4_r_v_b_1_80710 = net_80710;
  assign seg_20_17_sp4_r_v_b_30_80963 = seg_21_19_sp4_v_b_6_80963;
  assign seg_20_17_sp4_r_v_b_9_80718 = net_80718;
  assign seg_20_18_lutff_1_out_77468 = net_77468;
  assign seg_20_18_lutff_3_out_77470 = net_77470;
  assign seg_20_18_lutff_4_out_77471 = net_77471;
  assign seg_20_18_lutff_7_out_77474 = net_77474;
  assign seg_20_18_neigh_op_bnl_3_73904 = seg_19_17_ram_RDATA_12_73904;
  assign seg_20_18_neigh_op_bnl_5_73906 = seg_19_17_ram_RDATA_10_73906;
  assign seg_20_18_neigh_op_bnr_6_80938 = seg_21_17_lutff_6_out_80938;
  assign seg_20_18_neigh_op_lft_3_74027 = seg_19_18_ram_RDATA_4_74027;
  assign seg_20_18_neigh_op_lft_7_74031 = seg_19_18_ram_RDATA_0_74031;
  assign seg_20_18_neigh_op_top_6_77575 = seg_20_19_lutff_6_out_77575;
  assign seg_20_18_neigh_op_top_7_77576 = seg_20_19_lutff_7_out_77576;
  assign seg_20_18_sp4_h_l_43_66505 = seg_18_18_sp4_h_r_30_66505;
  assign seg_20_18_sp4_h_l_46_66500 = seg_17_18_sp4_h_r_22_66500;
  assign seg_20_18_sp4_r_v_b_27_81081 = net_81081;
  assign seg_20_19_lutff_6_out_77575 = net_77575;
  assign seg_20_19_lutff_7_out_77576 = net_77576;
  assign seg_20_19_sp4_h_r_45_70461 = seg_17_19_sp4_h_r_8_70461;
  assign seg_20_5_sp4_v_t_45_76408 = seg_20_7_sp4_v_b_32_76408;
  assign seg_20_6_lutff_2_out_76245 = net_76245;
  assign seg_20_6_lutff_5_out_76248 = net_76248;
  assign seg_20_6_lutff_7_out_76250 = net_76250;
  assign seg_20_6_neigh_op_rgt_5_79584 = seg_21_6_lutff_5_out_79584;
  assign seg_20_6_neigh_op_top_0_76345 = seg_20_7_lutff_0_out_76345;
  assign seg_20_6_sp4_h_r_26_72687 = seg_18_6_sp4_h_r_2_72687;
  assign seg_20_6_sp4_h_r_34_72685 = seg_18_6_sp4_h_r_10_72685;
  assign seg_20_6_sp4_h_r_4_79720 = net_79720;
  assign seg_20_6_sp4_r_v_b_33_79611 = net_79611;
  assign seg_20_6_sp4_v_t_43_76508 = seg_20_10_sp4_v_b_6_76508;
  assign seg_20_7_lutff_0_out_76345 = net_76345;
  assign seg_20_7_neigh_op_bnr_5_79584 = seg_21_6_lutff_5_out_79584;
  assign seg_20_7_sp4_h_r_16_76496 = net_76496;
  assign seg_20_7_sp4_r_v_b_1_79480 = net_79480;
  assign seg_20_7_sp4_r_v_b_33_79734 = net_79734;
  assign seg_20_7_sp4_v_b_26_76402 = seg_20_9_sp4_v_b_2_76402;
  assign seg_20_7_sp4_v_b_32_76408 = net_76408;
  assign seg_20_9_lutff_1_out_76550 = net_76550;
  assign seg_20_9_lutff_5_out_76554 = net_76554;
  assign seg_20_9_neigh_op_top_0_76651 = seg_20_10_lutff_0_out_76651;
  assign seg_20_9_neigh_op_top_3_76654 = seg_20_10_lutff_3_out_76654;
  assign seg_20_9_sp4_r_v_b_19_79856 = net_79856;
  assign seg_20_9_sp4_r_v_b_33_79980 = net_79980;
  assign seg_20_9_sp4_r_v_b_7_79732 = seg_21_6_sp4_v_b_42_79732;
  assign seg_20_9_sp4_v_b_2_76402 = net_76402;
  assign seg_21_10_lutff_0_out_80071 = net_80071;
  assign seg_21_10_lutff_1_out_80072 = net_80072;
  assign seg_21_10_lutff_4_out_80075 = net_80075;
  assign seg_21_10_neigh_op_bnl_5_76554 = seg_20_9_lutff_5_out_76554;
  assign seg_21_10_neigh_op_lft_0_76651 = seg_20_10_lutff_0_out_76651;
  assign seg_21_10_neigh_op_lft_3_76654 = seg_20_10_lutff_3_out_76654;
  assign seg_21_10_sp12_v_b_18_83666 = net_83666;
  assign seg_21_10_sp4_h_r_10_84039 = net_84039;
  assign seg_21_10_sp4_h_r_13_80206 = seg_20_10_sp4_h_r_0_80206;
  assign seg_21_10_sp4_h_r_18_80215 = net_80215;
  assign seg_21_10_sp4_h_r_24_76795 = net_76795;
  assign seg_21_10_sp4_h_r_2_84041 = net_84041;
  assign seg_21_10_sp4_h_r_34_76797 = net_76797;
  assign seg_21_10_sp4_h_r_8_84047 = net_84047;
  assign seg_21_10_sp4_r_v_b_25_83926 = net_83926;
  assign seg_21_10_sp4_v_b_18_79978 = net_79978;
  assign seg_21_10_sp4_v_b_24_80096 = net_80096;
  assign seg_21_10_sp4_v_b_34_80106 = net_80106;
  assign seg_21_10_sp4_v_b_40_80222 = net_80222;
  assign seg_21_10_sp4_v_b_6_79856 = seg_20_9_sp4_r_v_b_19_79856;
  assign seg_21_11_sp4_v_b_2_79975 = seg_20_10_sp4_r_v_b_15_79975;
  assign seg_21_11_sp4_v_b_7_79978 = seg_21_10_sp4_v_b_18_79978;
  assign seg_21_11_sp4_v_t_36_80464 = seg_21_14_sp4_v_b_12_80464;
  assign seg_21_12_lutff_2_out_80319 = net_80319;
  assign seg_21_12_lutff_7_out_80324 = net_80324;
  assign seg_21_12_neigh_op_lft_0_76855 = seg_20_12_lutff_0_out_76855;
  assign seg_21_12_neigh_op_lft_7_76862 = seg_20_12_lutff_7_out_76862;
  assign seg_21_12_sp4_v_b_0_80096 = seg_21_10_sp4_v_b_24_80096;
  assign seg_21_12_sp4_v_b_10_80106 = seg_21_10_sp4_v_b_34_80106;
  assign seg_21_12_sp4_v_b_16_80222 = seg_21_10_sp4_v_b_40_80222;
  assign seg_21_12_sp4_v_b_1_80095 = seg_21_9_sp4_v_b_36_80095;
  assign seg_21_12_sp4_v_b_23_80229 = seg_20_10_sp4_r_v_b_47_80229;
  assign seg_21_12_sp4_v_b_42_80470 = net_80470;
  assign seg_21_12_sp4_v_b_7_80101 = seg_20_10_sp4_r_v_b_31_80101;
  assign seg_21_13_lutff_1_out_80441 = net_80441;
  assign seg_21_13_lutff_2_out_80442 = net_80442;
  assign seg_21_13_lutff_6_out_80446 = net_80446;
  assign seg_21_13_lutff_7_out_80447 = net_80447;
  assign seg_21_13_neigh_op_bot_2_80319 = seg_21_12_lutff_2_out_80319;
  assign seg_21_13_neigh_op_lft_4_76961 = seg_20_13_lutff_4_out_76961;
  assign seg_21_13_neigh_op_rgt_2_84273 = seg_22_13_lutff_2_out_84273;
  assign seg_21_13_sp4_h_l_42_69722 = seg_20_13_sp4_h_r_42_69722;
  assign seg_21_13_sp4_h_l_46_69716 = seg_18_13_sp4_h_r_22_69716;
  assign seg_21_13_sp4_h_r_24_77101 = seg_19_13_sp4_h_r_0_77101;
  assign seg_21_13_sp4_h_r_31_77110 = seg_22_13_sp4_h_r_42_77110;
  assign seg_21_13_sp4_h_r_37_73544 = seg_18_13_sp4_h_r_0_73544;
  assign seg_21_13_sp4_h_r_45_73554 = seg_18_13_sp4_h_r_8_73554;
  assign seg_21_13_sp4_r_v_b_41_84423 = net_84423;
  assign seg_21_13_sp4_v_b_10_80229 = seg_20_10_sp4_r_v_b_47_80229;
  assign seg_21_13_sp4_v_b_32_80473 = net_80473;
  assign seg_21_13_sp4_v_b_38_80589 = net_80589;
  assign seg_21_13_sp4_v_b_5_80222 = seg_21_10_sp4_v_b_40_80222;
  assign seg_21_14_lutff_1_out_80564 = net_80564;
  assign seg_21_14_lutff_2_out_80565 = net_80565;
  assign seg_21_14_lutff_3_out_80566 = net_80566;
  assign seg_21_14_lutff_4_out_80567 = net_80567;
  assign seg_21_14_lutff_5_out_80568 = net_80568;
  assign seg_21_14_lutff_7_out_80570 = net_80570;
  assign seg_21_14_neigh_op_bnl_0_76957 = seg_20_13_lutff_0_out_76957;
  assign seg_21_14_neigh_op_bot_2_80442 = seg_21_13_lutff_2_out_80442;
  assign seg_21_14_neigh_op_lft_3_77062 = seg_20_14_lutff_3_out_77062;
  assign seg_21_14_neigh_op_lft_7_77066 = seg_20_14_lutff_7_out_77066;
  assign seg_21_14_neigh_op_top_0_80686 = seg_21_15_lutff_0_out_80686;
  assign seg_21_14_neigh_op_top_1_80687 = seg_21_15_lutff_1_out_80687;
  assign seg_21_14_neigh_op_top_5_80691 = seg_21_15_lutff_5_out_80691;
  assign seg_21_14_neigh_op_top_7_80693 = seg_21_15_lutff_7_out_80693;
  assign seg_21_14_sp12_v_b_11_83667 = seg_21_9_sp12_v_b_20_83667;
  assign seg_21_14_sp4_v_b_12_80464 = net_80464;
  assign seg_21_14_sp4_v_b_18_80470 = seg_21_12_sp4_v_b_42_80470;
  assign seg_21_14_sp4_v_b_32_80596 = net_80596;
  assign seg_21_14_sp4_v_b_36_80710 = seg_20_17_sp4_r_v_b_1_80710;
  assign seg_21_14_sp4_v_b_44_80718 = seg_20_17_sp4_r_v_b_9_80718;
  assign seg_21_14_sp4_v_t_36_80833 = seg_21_17_sp4_v_b_12_80833;
  assign seg_21_14_sp4_v_t_47_80844 = seg_21_18_sp4_v_b_10_80844;
  assign seg_21_15_lutff_0_out_80686 = net_80686;
  assign seg_21_15_lutff_1_out_80687 = net_80687;
  assign seg_21_15_lutff_2_out_80688 = net_80688;
  assign seg_21_15_lutff_3_out_80689 = net_80689;
  assign seg_21_15_lutff_4_out_80690 = net_80690;
  assign seg_21_15_lutff_5_out_80691 = net_80691;
  assign seg_21_15_lutff_6_out_80692 = net_80692;
  assign seg_21_15_lutff_7_out_80693 = net_80693;
  assign seg_21_15_neigh_op_lft_0_77161 = seg_20_15_lutff_0_out_77161;
  assign seg_21_15_neigh_op_lft_2_77163 = seg_20_15_lutff_2_out_77163;
  assign seg_21_15_neigh_op_lft_3_77164 = seg_20_15_lutff_3_out_77164;
  assign seg_21_15_neigh_op_lft_5_77166 = seg_20_15_lutff_5_out_77166;
  assign seg_21_15_neigh_op_tnr_7_84647 = seg_22_16_lutff_7_out_84647;
  assign seg_21_15_neigh_op_top_3_80812 = seg_21_16_lutff_3_out_80812;
  assign seg_21_15_sp4_h_l_43_69967 = seg_17_15_sp4_h_r_6_69967;
  assign seg_21_15_sp4_r_v_b_17_84423 = seg_21_13_sp4_r_v_b_41_84423;
  assign seg_21_15_sp4_v_b_14_80589 = seg_21_13_sp4_v_b_38_80589;
  assign seg_21_15_sp4_v_b_21_80596 = seg_21_14_sp4_v_b_32_80596;
  assign seg_21_15_sp4_v_b_41_80838 = seg_21_18_sp4_v_b_4_80838;
  assign seg_21_15_sp4_v_b_8_80473 = seg_21_13_sp4_v_b_32_80473;
  assign seg_21_15_sp4_v_t_38_80958 = seg_21_18_sp4_v_b_14_80958;
  assign seg_21_16_lutff_3_out_80812 = net_80812;
  assign seg_21_16_lutff_4_out_80813 = net_80813;
  assign seg_21_16_lutff_6_out_80815 = net_80815;
  assign seg_21_16_neigh_op_tnl_1_77366 = seg_20_17_lutff_1_out_77366;
  assign seg_21_16_neigh_op_top_5_80937 = seg_21_17_lutff_5_out_80937;
  assign seg_21_16_sp4_h_l_39_70086 = seg_19_16_sp4_h_r_26_70086;
  assign seg_21_16_sp4_h_l_44_70093 = seg_18_16_sp4_h_r_20_70093;
  assign seg_21_16_sp4_h_r_24_77407 = net_77407;
  assign seg_21_16_sp4_v_t_38_81081 = seg_20_18_sp4_r_v_b_27_81081;
  assign seg_21_17_lutff_0_out_80932 = net_80932;
  assign seg_21_17_lutff_1_out_80933 = net_80933;
  assign seg_21_17_lutff_2_out_80934 = net_80934;
  assign seg_21_17_lutff_3_out_80935 = net_80935;
  assign seg_21_17_lutff_4_out_80936 = net_80936;
  assign seg_21_17_lutff_5_out_80937 = net_80937;
  assign seg_21_17_lutff_6_out_80938 = net_80938;
  assign seg_21_17_lutff_7_out_80939 = net_80939;
  assign seg_21_17_neigh_op_bnl_1_77264 = seg_20_16_lutff_1_out_77264;
  assign seg_21_17_neigh_op_bnl_2_77265 = seg_20_16_lutff_2_out_77265;
  assign seg_21_17_neigh_op_bnl_3_77266 = seg_20_16_lutff_3_out_77266;
  assign seg_21_17_neigh_op_bnl_6_77269 = seg_20_16_lutff_6_out_77269;
  assign seg_21_17_neigh_op_bnl_7_77270 = seg_20_16_lutff_7_out_77270;
  assign seg_21_17_neigh_op_bot_4_80813 = seg_21_16_lutff_4_out_80813;
  assign seg_21_17_neigh_op_lft_2_77367 = seg_20_17_lutff_2_out_77367;
  assign seg_21_17_neigh_op_rgt_2_84765 = seg_22_17_lutff_2_out_84765;
  assign seg_21_17_neigh_op_rgt_5_84768 = seg_22_17_lutff_5_out_84768;
  assign seg_21_17_neigh_op_rgt_6_84769 = seg_22_17_lutff_6_out_84769;
  assign seg_21_17_sp4_h_l_36_70206 = seg_18_17_sp4_h_r_12_70206;
  assign seg_21_17_sp4_h_r_11_84901 = seg_22_17_sp4_h_r_22_84901;
  assign seg_21_17_sp4_h_r_12_81068 = net_81068;
  assign seg_21_17_sp4_h_r_1_84899 = seg_22_17_sp4_h_r_12_84899;
  assign seg_21_17_sp4_h_r_37_74036 = seg_18_17_sp4_h_r_0_74036;
  assign seg_21_17_sp4_h_r_3_84903 = seg_22_17_sp4_h_r_14_84903;
  assign seg_21_17_sp4_h_r_41_74042 = seg_18_17_sp4_h_r_4_74042;
  assign seg_21_17_sp4_h_r_44_74047 = net_74047;
  assign seg_21_17_sp4_h_r_7_84907 = seg_22_17_sp4_h_r_18_84907;
  assign seg_21_17_sp4_r_v_b_12_84664 = seg_22_15_sp4_v_b_36_84664;
  assign seg_21_17_sp4_r_v_b_13_84665 = net_84665;
  assign seg_21_17_sp4_v_b_12_80833 = net_80833;
  assign seg_21_18_lutff_1_out_81056 = net_81056;
  assign seg_21_18_lutff_3_out_81058 = net_81058;
  assign seg_21_18_lutff_4_out_81059 = net_81059;
  assign seg_21_18_lutff_6_out_81061 = net_81061;
  assign seg_21_18_neigh_op_lft_1_77468 = seg_20_18_lutff_1_out_77468;
  assign seg_21_18_neigh_op_lft_3_77470 = seg_20_18_lutff_3_out_77470;
  assign seg_21_18_neigh_op_lft_4_77471 = seg_20_18_lutff_4_out_77471;
  assign seg_21_18_neigh_op_top_2_81180 = seg_21_19_lutff_2_out_81180;
  assign seg_21_18_sp12_h_r_8_70324 = net_70324;
  assign seg_21_18_sp12_v_b_2_83666 = seg_21_10_sp12_v_b_18_83666;
  assign seg_21_18_sp4_h_l_36_70329 = seg_18_18_sp4_h_r_12_70329;
  assign seg_21_18_sp4_h_r_41_74165 = seg_18_18_sp4_h_r_4_74165;
  assign seg_21_18_sp4_v_b_10_80844 = net_80844;
  assign seg_21_18_sp4_v_b_14_80958 = net_80958;
  assign seg_21_18_sp4_v_b_1_80833 = seg_21_17_sp4_v_b_12_80833;
  assign seg_21_18_sp4_v_b_3_80835 = seg_20_16_sp4_r_v_b_27_80835;
  assign seg_21_18_sp4_v_b_4_80838 = net_80838;
  assign seg_21_18_sp4_v_b_7_80839 = seg_20_16_sp4_r_v_b_31_80839;
  assign seg_21_19_lutff_2_out_81180 = net_81180;
  assign seg_21_19_sp4_v_b_6_80963 = net_80963;
  assign seg_21_5_sp4_v_t_44_79734 = seg_20_7_sp4_r_v_b_33_79734;
  assign seg_21_6_lutff_5_out_79584 = net_79584;
  assign seg_21_6_neigh_op_lft_5_76248 = seg_20_6_lutff_5_out_76248;
  assign seg_21_6_neigh_op_lft_7_76250 = seg_20_6_lutff_7_out_76250;
  assign seg_21_6_sp12_v_b_10_82776 = net_82776;
  assign seg_21_6_sp4_h_r_10_83547 = net_83547;
  assign seg_21_6_sp4_h_r_26_76391 = net_76391;
  assign seg_21_6_sp4_h_r_42_72692 = net_72692;
  assign seg_21_6_sp4_r_v_b_11_83198 = net_83198;
  assign seg_21_6_sp4_r_v_b_43_83564 = net_83564;
  assign seg_21_6_sp4_r_v_b_7_83194 = net_83194;
  assign seg_21_6_sp4_v_b_10_79368 = net_79368;
  assign seg_21_6_sp4_v_b_42_79732 = net_79732;
  assign seg_21_7_sp4_v_b_1_79480 = seg_20_7_sp4_r_v_b_1_79480;
  assign seg_21_9_lutff_0_out_79948 = net_79948;
  assign seg_21_9_lutff_2_out_79950 = net_79950;
  assign seg_21_9_neigh_op_lft_5_76554 = seg_20_9_lutff_5_out_76554;
  assign seg_21_9_sp12_v_b_20_83667 = net_83667;
  assign seg_21_9_sp12_v_b_5_82776 = seg_21_6_sp12_v_b_10_82776;
  assign seg_21_9_sp4_h_r_0_83914 = net_83914;
  assign seg_21_9_sp4_h_r_20_80094 = net_80094;
  assign seg_21_9_sp4_h_r_28_76699 = net_76699;
  assign seg_21_9_sp4_v_b_36_80095 = net_80095;
  assign seg_21_9_sp4_v_b_7_79732 = seg_21_6_sp4_v_b_42_79732;
  assign seg_22_10_sp4_h_l_43_73183 = seg_18_10_sp4_h_r_6_73183;
  assign seg_22_12_sp4_v_b_1_83926 = seg_21_10_sp4_r_v_b_25_83926;
  assign seg_22_13_lutff_2_out_84273 = net_84273;
  assign seg_22_13_sp4_h_r_42_77110 = net_77110;
  assign seg_22_13_sp4_v_t_43_84548 = seg_22_17_sp4_v_b_6_84548;
  assign seg_22_13_sp4_v_t_45_84550 = seg_22_17_sp4_v_b_8_84550;
  assign seg_22_14_neigh_op_top_4_84521 = seg_22_15_lutff_4_out_84521;
  assign seg_22_14_sp4_h_l_40_73674 = seg_19_14_sp4_h_r_16_73674;
  assign seg_22_14_sp4_h_r_38_77208 = net_77208;
  assign seg_22_14_sp4_v_t_37_84665 = seg_21_17_sp4_r_v_b_13_84665;
  assign seg_22_15_lutff_4_out_84521 = net_84521;
  assign seg_22_15_sp4_h_l_38_73795 = seg_19_15_sp4_h_r_14_73795;
  assign seg_22_15_sp4_r_v_b_37_88496 = net_88496;
  assign seg_22_15_sp4_v_b_36_84664 = net_84664;
  assign seg_22_15_sp4_v_b_38_84666 = seg_22_17_sp4_v_b_14_84666;
  assign seg_22_15_sp4_v_t_41_84792 = seg_22_17_sp4_v_b_28_84792;
  assign seg_22_15_sp4_v_t_47_84798 = seg_22_17_sp4_v_b_34_84798;
  assign seg_22_16_lutff_7_out_84647 = net_84647;
  assign seg_22_16_neigh_op_tnl_6_80938 = seg_21_17_lutff_6_out_80938;
  assign seg_22_17_lutff_2_out_84765 = net_84765;
  assign seg_22_17_lutff_5_out_84768 = net_84768;
  assign seg_22_17_lutff_6_out_84769 = net_84769;
  assign seg_22_17_neigh_op_lft_3_80935 = seg_21_17_lutff_3_out_80935;
  assign seg_22_17_neigh_op_lft_4_80936 = seg_21_17_lutff_4_out_80936;
  assign seg_22_17_neigh_op_lft_5_80937 = seg_21_17_lutff_5_out_80937;
  assign seg_22_17_neigh_op_lft_7_80939 = seg_21_17_lutff_7_out_80939;
  assign seg_22_17_sp4_h_l_37_74036 = seg_18_17_sp4_h_r_0_74036;
  assign seg_22_17_sp4_h_l_41_74042 = seg_18_17_sp4_h_r_4_74042;
  assign seg_22_17_sp4_h_l_47_74038 = seg_18_17_sp4_h_r_10_74038;
  assign seg_22_17_sp4_h_r_12_84899 = net_84899;
  assign seg_22_17_sp4_h_r_14_84903 = net_84903;
  assign seg_22_17_sp4_h_r_18_84907 = net_84907;
  assign seg_22_17_sp4_h_r_22_84901 = net_84901;
  assign seg_22_17_sp4_h_r_36_77510 = net_77510;
  assign seg_22_17_sp4_h_r_38_77514 = net_77514;
  assign seg_22_17_sp4_h_r_40_77516 = net_77516;
  assign seg_22_17_sp4_h_r_42_77518 = net_77518;
  assign seg_22_17_sp4_h_r_46_77512 = net_77512;
  assign seg_22_17_sp4_h_r_8_88739 = net_88739;
  assign seg_22_17_sp4_r_v_b_11_88382 = net_88382;
  assign seg_22_17_sp4_r_v_b_13_88496 = seg_22_15_sp4_r_v_b_37_88496;
  assign seg_22_17_sp4_r_v_b_3_88374 = net_88374;
  assign seg_22_17_sp4_r_v_b_5_88376 = net_88376;
  assign seg_22_17_sp4_v_b_14_84666 = net_84666;
  assign seg_22_17_sp4_v_b_28_84792 = net_84792;
  assign seg_22_17_sp4_v_b_2_84544 = net_84544;
  assign seg_22_17_sp4_v_b_34_84798 = net_84798;
  assign seg_22_17_sp4_v_b_6_84548 = net_84548;
  assign seg_22_17_sp4_v_b_8_84550 = net_84550;
  assign seg_22_2_sp4_v_t_42_83194 = seg_21_6_sp4_r_v_b_7_83194;
  assign seg_22_6_sp4_h_l_39_72687 = seg_18_6_sp4_h_r_2_72687;
  assign seg_22_6_sp4_v_b_11_83198 = seg_21_6_sp4_r_v_b_11_83198;
  assign seg_22_9_lutff_1_out_83780 = net_83780;
  assign seg_22_9_sp4_v_b_6_83564 = seg_21_6_sp4_r_v_b_43_83564;
  assign seg_23_13_sp4_v_t_38_88374 = seg_22_17_sp4_r_v_b_3_88374;
  assign seg_23_13_sp4_v_t_40_88376 = seg_22_17_sp4_r_v_b_5_88376;
  assign seg_23_13_sp4_v_t_46_88382 = seg_22_17_sp4_r_v_b_11_88382;
  assign seg_23_17_sp4_h_l_37_77509 = seg_19_17_sp4_h_r_0_77509;
  assign seg_23_6_sp4_v_t_38_87513 = seg_23_9_sp4_v_b_14_87513;
  assign seg_23_9_lutff_2_out_87612 = net_87612;
  assign seg_23_9_neigh_op_lft_1_83780 = seg_22_9_lutff_1_out_83780;
  assign seg_23_9_sp4_h_l_41_76699 = seg_21_9_sp4_h_r_28_76699;
  assign seg_23_9_sp4_h_r_24_83914 = seg_21_9_sp4_h_r_0_83914;
  assign seg_23_9_sp4_v_b_14_87513 = net_87513;
  assign seg_24_9_sp4_h_l_44_80094 = seg_21_9_sp4_h_r_20_80094;
  assign seg_2_19_neigh_op_rgt_4_13488 = seg_3_19_lutff_4_out_13488;
  assign seg_2_19_neigh_op_rgt_5_13489 = seg_3_19_lutff_5_out_13489;
  assign seg_2_19_neigh_op_rgt_6_13490 = seg_3_19_lutff_6_out_13490;
  assign seg_2_19_neigh_op_tnr_2_13609 = seg_3_20_lutff_2_out_13609;
  assign seg_2_19_sp4_h_r_0_13619 = net_13619;
  assign seg_2_8_lutff_2_out_7745 = net_7745;
  assign seg_2_8_lutff_3_out_7746 = net_7746;
  assign seg_2_8_lutff_4_out_7747 = net_7747;
  assign seg_2_8_lutff_5_out_7748 = net_7748;
  assign seg_2_8_lutff_6_out_7749 = net_7749;
  assign seg_2_8_neigh_op_bnr_7_12015 = seg_3_7_lutff_7_out_12015;
  assign seg_2_8_neigh_op_rgt_4_12135 = seg_3_8_lutff_4_out_12135;
  assign seg_2_8_sp4_h_r_46_1816 = net_1816;
  assign seg_2_8_sp4_r_v_b_15_12035 = net_12035;
  assign seg_3_13_lutff_2_out_12748 = net_12748;
  assign seg_3_13_lutff_3_out_12749 = net_12749;
  assign seg_3_13_lutff_4_out_12750 = net_12750;
  assign seg_3_13_lutff_5_out_12751 = net_12751;
  assign seg_3_13_lutff_6_out_12752 = net_12752;
  assign seg_3_13_neigh_op_rgt_5_16582 = seg_4_13_lutff_5_out_16582;
  assign seg_3_13_neigh_op_top_2_12871 = seg_3_14_lutff_2_out_12871;
  assign seg_3_13_sp12_v_b_14_16095 = net_16095;
  assign seg_3_13_sp4_h_r_14_12886 = net_12886;
  assign seg_3_13_sp4_h_r_46_2864 = net_2864;
  assign seg_3_14_lutff_2_out_12871 = net_12871;
  assign seg_3_14_sp12_v_b_13_16095 = seg_3_13_sp12_v_b_14_16095;
  assign seg_3_18_lutff_2_out_13363 = net_13363;
  assign seg_3_18_lutff_3_out_13364 = net_13364;
  assign seg_3_18_lutff_4_out_13365 = net_13365;
  assign seg_3_18_lutff_5_out_13366 = net_13366;
  assign seg_3_18_lutff_6_out_13367 = net_13367;
  assign seg_3_18_lutff_7_out_13368 = net_13368;
  assign seg_3_18_neigh_op_bnr_1_17070 = seg_4_17_lutff_1_out_17070;
  assign seg_3_18_neigh_op_rgt_7_17199 = seg_4_18_lutff_7_out_17199;
  assign seg_3_19_lutff_0_out_13484 = net_13484;
  assign seg_3_19_lutff_1_out_13485 = net_13485;
  assign seg_3_19_lutff_2_out_13486 = net_13486;
  assign seg_3_19_lutff_3_out_13487 = net_13487;
  assign seg_3_19_lutff_4_out_13488 = net_13488;
  assign seg_3_19_lutff_5_out_13489 = net_13489;
  assign seg_3_19_lutff_6_out_13490 = net_13490;
  assign seg_3_19_lutff_7_out_13491 = net_13491;
  assign seg_3_20_lutff_0_out_13607 = net_13607;
  assign seg_3_20_lutff_1_out_13608 = net_13608;
  assign seg_3_20_lutff_2_out_13609 = net_13609;
  assign seg_3_20_lutff_3_out_13610 = net_13610;
  assign seg_3_20_lutff_4_out_13611 = net_13611;
  assign seg_3_20_lutff_5_out_13612 = net_13612;
  assign seg_3_20_lutff_6_out_13613 = net_13613;
  assign seg_3_20_lutff_7_out_13614 = net_13614;
  assign seg_3_5_sp4_v_t_39_12035 = seg_2_8_sp4_r_v_b_15_12035;
  assign seg_3_7_lutff_7_out_12015 = net_12015;
  assign seg_3_7_sp4_v_b_30_12039 = net_12039;
  assign seg_3_8_lutff_4_out_12135 = net_12135;
  assign seg_3_8_sp4_h_l_46_1816 = seg_2_8_sp4_h_r_46_1816;
  assign seg_3_8_sp4_v_b_19_12039 = seg_3_7_sp4_v_b_30_12039;
  assign seg_4_12_lutff_2_out_16456 = net_16456;
  assign seg_4_12_sp4_h_r_4_20426 = net_20426;
  assign seg_4_13_lutff_5_out_16582 = net_16582;
  assign seg_4_13_sp4_h_l_46_2864 = seg_3_13_sp4_h_r_46_2864;
  assign seg_4_13_sp4_v_b_10_16366 = net_16366;
  assign seg_4_17_lutff_1_out_17070 = net_17070;
  assign seg_4_17_sp4_v_b_27_17095 = seg_4_18_sp4_v_b_14_17095;
  assign seg_4_18_lutff_0_out_17192 = net_17192;
  assign seg_4_18_lutff_6_out_17198 = net_17198;
  assign seg_4_18_lutff_7_out_17199 = net_17199;
  assign seg_4_18_neigh_op_bot_1_17070 = seg_4_17_lutff_1_out_17070;
  assign seg_4_18_neigh_op_lft_2_13363 = seg_3_18_lutff_2_out_13363;
  assign seg_4_18_neigh_op_lft_3_13364 = seg_3_18_lutff_3_out_13364;
  assign seg_4_18_neigh_op_lft_4_13365 = seg_3_18_lutff_4_out_13365;
  assign seg_4_18_neigh_op_lft_5_13366 = seg_3_18_lutff_5_out_13366;
  assign seg_4_18_neigh_op_lft_6_13367 = seg_3_18_lutff_6_out_13367;
  assign seg_4_18_neigh_op_tnl_1_13485 = seg_3_19_lutff_1_out_13485;
  assign seg_4_18_neigh_op_top_1_17316 = seg_4_19_lutff_1_out_17316;
  assign seg_4_18_sp4_h_r_4_21164 = net_21164;
  assign seg_4_18_sp4_r_v_b_21_20933 = net_20933;
  assign seg_4_18_sp4_r_v_b_37_21171 = net_21171;
  assign seg_4_18_sp4_r_v_b_5_20805 = net_20805;
  assign seg_4_18_sp4_v_b_14_17095 = net_17095;
  assign seg_4_19_lutff_1_out_17316 = net_17316;
  assign seg_4_19_lutff_2_out_17317 = net_17317;
  assign seg_4_19_lutff_4_out_17319 = net_17319;
  assign seg_4_19_neigh_op_bnl_7_13368 = seg_3_18_lutff_7_out_13368;
  assign seg_4_19_neigh_op_lft_0_13484 = seg_3_19_lutff_0_out_13484;
  assign seg_4_19_neigh_op_lft_2_13486 = seg_3_19_lutff_2_out_13486;
  assign seg_4_19_neigh_op_lft_3_13487 = seg_3_19_lutff_3_out_13487;
  assign seg_4_19_neigh_op_lft_7_13491 = seg_3_19_lutff_7_out_13491;
  assign seg_4_19_neigh_op_tnl_0_13607 = seg_3_20_lutff_0_out_13607;
  assign seg_4_19_neigh_op_tnl_5_13612 = seg_3_20_lutff_5_out_13612;
  assign seg_4_19_neigh_op_tnl_7_13614 = seg_3_20_lutff_7_out_13614;
  assign seg_4_19_neigh_op_top_1_17439 = seg_4_20_lutff_1_out_17439;
  assign seg_4_19_sp4_h_r_24_13619 = seg_2_19_sp4_h_r_0_13619;
  assign seg_4_20_lutff_1_out_17439 = net_17439;
  assign seg_4_20_neigh_op_lft_1_13608 = seg_3_20_lutff_1_out_13608;
  assign seg_4_20_neigh_op_lft_3_13610 = seg_3_20_lutff_3_out_13610;
  assign seg_4_20_neigh_op_lft_4_13611 = seg_3_20_lutff_4_out_13611;
  assign seg_4_20_neigh_op_lft_6_13613 = seg_3_20_lutff_6_out_13613;
  assign seg_5_12_lutff_2_out_20287 = net_20287;
  assign seg_5_12_neigh_op_lft_2_16456 = seg_4_12_lutff_2_out_16456;
  assign seg_5_12_sp4_h_r_4_24257 = net_24257;
  assign seg_5_14_sp4_v_t_40_20805 = seg_4_18_sp4_r_v_b_5_20805;
  assign seg_5_17_sp4_v_t_37_21171 = seg_4_18_sp4_r_v_b_37_21171;
  assign seg_5_19_sp4_v_b_8_20933 = seg_4_18_sp4_r_v_b_21_20933;
  assign seg_5_20_sp12_h_r_3_21400 = seg_10_20_sp12_h_r_12_21400;
  assign seg_5_20_sp4_h_r_4_25241 = net_25241;
  assign seg_5_5_sp4_h_r_0_23390 = net_23390;
  assign seg_5_5_sp4_r_v_b_17_23161 = net_23161;
  assign seg_6_0_span12_vert_18_26571 = net_26571;
  assign seg_6_0_span4_vert_32_22900 = net_22900;
  assign seg_6_10_sp12_v_b_1_26571 = seg_6_0_span12_vert_18_26571;
  assign seg_6_13_sp4_h_l_38_12886 = seg_3_13_sp4_h_r_14_12886;
  assign seg_6_2_sp4_h_r_2_26813 = seg_8_2_sp4_h_r_26_26813;
  assign seg_6_2_sp4_v_t_41_23161 = seg_5_5_sp4_r_v_b_17_23161;
  assign seg_6_3_sp4_v_b_8_22900 = seg_6_0_span4_vert_32_22900;
  assign seg_6_4_sp4_h_r_10_27015 = seg_8_4_sp4_h_r_34_27015;
  assign seg_7_0_span4_vert_16_26691 = net_26691;
  assign seg_7_10_sp4_h_r_3_31041 = seg_8_10_sp4_h_r_14_31041;
  assign seg_7_12_lutff_2_out_27687 = net_27687;
  assign seg_7_12_lutff_3_out_27688 = net_27688;
  assign seg_7_12_sp4_h_r_10_31284 = net_31284;
  assign seg_7_12_sp4_h_r_28_24257 = seg_5_12_sp4_h_r_4_24257;
  assign seg_7_12_sp4_h_r_41_20426 = seg_4_12_sp4_h_r_4_20426;
  assign seg_7_1_neigh_op_tnr_3_29884 = seg_8_2_lutff_3_out_29884;
  assign seg_7_1_neigh_op_tnr_7_29888 = seg_8_2_lutff_7_out_29888;
  assign seg_7_2_sp4_v_b_5_26691 = seg_7_0_span4_vert_16_26691;
  assign seg_7_4_sp4_h_r_7_30307 = seg_8_4_sp4_h_r_18_30307;
  assign seg_8_0_span4_vert_37_29936 = seg_8_2_sp4_v_b_24_29936;
  assign seg_8_10_lutff_2_out_30903 = net_30903;
  assign seg_8_10_lutff_3_out_30904 = net_30904;
  assign seg_8_10_lutff_4_out_30905 = net_30905;
  assign seg_8_10_lutff_5_out_30906 = net_30906;
  assign seg_8_10_lutff_6_out_30907 = net_30907;
  assign seg_8_10_neigh_op_top_5_31029 = seg_8_11_lutff_5_out_31029;
  assign seg_8_10_sp12_v_b_14_34250 = net_34250;
  assign seg_8_10_sp4_h_r_14_31041 = net_31041;
  assign seg_8_10_sp4_h_r_30_27633 = net_27633;
  assign seg_8_10_sp4_h_r_46_24008 = net_24008;
  assign seg_8_10_sp4_v_b_26_30928 = seg_8_12_sp4_v_b_2_30928;
  assign seg_8_11_lutff_5_out_31029 = net_31029;
  assign seg_8_11_sp12_v_b_13_34250 = seg_8_10_sp12_v_b_14_34250;
  assign seg_8_12_lutff_1_out_31148 = net_31148;
  assign seg_8_12_sp12_v_b_2_33722 = seg_8_4_sp12_v_b_18_33722;
  assign seg_8_12_sp4_h_r_2_35117 = net_35117;
  assign seg_8_12_sp4_v_b_2_30928 = net_30928;
  assign seg_8_13_sp12_v_b_1_33722 = seg_8_4_sp12_v_b_18_33722;
  assign seg_8_17_sp4_h_r_26_28343 = net_28343;
  assign seg_8_17_sp4_r_v_b_43_35747 = net_35747;
  assign seg_8_18_sp4_h_l_41_21164 = seg_4_18_sp4_h_r_4_21164;
  assign seg_8_23_lutff_5_out_32505 = net_32505;
  assign seg_8_23_sp4_v_b_26_32527 = net_32527;
  assign seg_8_23_sp4_v_t_41_32775 = seg_8_25_sp4_v_b_28_32775;
  assign seg_8_24_lutff_6_out_32629 = net_32629;
  assign seg_8_24_sp4_v_t_44_32901 = seg_8_25_sp4_v_b_44_32901;
  assign seg_8_25_lutff_2_out_32748 = net_32748;
  assign seg_8_25_lutff_3_out_32749 = net_32749;
  assign seg_8_25_lutff_4_out_32750 = net_32750;
  assign seg_8_25_lutff_5_out_32751 = net_32751;
  assign seg_8_25_lutff_7_out_32753 = net_32753;
  assign seg_8_25_neigh_op_bot_6_32629 = seg_8_24_lutff_6_out_32629;
  assign seg_8_25_sp4_h_r_12_32882 = net_32882;
  assign seg_8_25_sp4_r_v_b_29_36605 = net_36605;
  assign seg_8_25_sp4_v_b_28_32775 = net_32775;
  assign seg_8_25_sp4_v_b_2_32527 = seg_8_23_sp4_v_b_26_32527;
  assign seg_8_25_sp4_v_b_44_32901 = net_32901;
  assign seg_8_2_lutff_1_out_29882 = net_29882;
  assign seg_8_2_lutff_2_out_29883 = net_29883;
  assign seg_8_2_lutff_3_out_29884 = net_29884;
  assign seg_8_2_lutff_6_out_29887 = net_29887;
  assign seg_8_2_lutff_7_out_29888 = net_29888;
  assign seg_8_2_neigh_op_rgt_0_33712 = seg_9_2_lutff_0_out_33712;
  assign seg_8_2_neigh_op_tnr_1_33872 = seg_9_3_lutff_1_out_33872;
  assign seg_8_2_neigh_op_tnr_2_33873 = seg_9_3_lutff_2_out_33873;
  assign seg_8_2_neigh_op_tnr_4_33875 = seg_9_3_lutff_4_out_33875;
  assign seg_8_2_neigh_op_top_5_30045 = seg_8_3_lutff_5_out_30045;
  assign seg_8_2_sp4_h_r_26_26813 = net_26813;
  assign seg_8_2_sp4_v_b_24_29936 = net_29936;
  assign seg_8_30_sp4_v_t_36_37347 = seg_8_31_span4_vert_36_37347;
  assign seg_8_31_io_1_D_IN_0_33486 = net_33486;
  assign seg_8_31_logic_op_bnr_7_37199 = seg_9_30_lutff_7_out_37199;
  assign seg_8_31_span4_horz_r_6_33556 = net_33556;
  assign seg_8_31_span4_vert_36_37347 = net_37347;
  assign seg_8_3_lutff_4_out_30044 = net_30044;
  assign seg_8_3_lutff_5_out_30045 = net_30045;
  assign seg_8_3_lutff_6_out_30046 = net_30046;
  assign seg_8_3_neigh_op_rgt_1_33872 = seg_9_3_lutff_1_out_33872;
  assign seg_8_3_neigh_op_rgt_2_33873 = seg_9_3_lutff_2_out_33873;
  assign seg_8_3_neigh_op_rgt_4_33875 = seg_9_3_lutff_4_out_33875;
  assign seg_8_3_sp4_h_r_18_30184 = net_30184;
  assign seg_8_3_sp4_h_r_30_26919 = net_26919;
  assign seg_8_3_sp4_r_v_b_19_33774 = net_33774;
  assign seg_8_4_lutff_1_out_30164 = net_30164;
  assign seg_8_4_sp12_v_b_18_33722 = net_33722;
  assign seg_8_4_sp4_h_r_18_30307 = net_30307;
  assign seg_8_4_sp4_h_r_2_34133 = net_34133;
  assign seg_8_4_sp4_h_r_34_27015 = net_27015;
  assign seg_8_4_sp4_r_v_b_35_34028 = net_34028;
  assign seg_8_4_sp4_r_v_b_3_33768 = net_33768;
  assign seg_8_4_sp4_v_b_34_30198 = net_30198;
  assign seg_8_6_sp4_v_b_10_30198 = seg_8_4_sp4_v_b_34_30198;
  assign seg_9_10_lutff_1_out_34733 = net_34733;
  assign seg_9_10_lutff_2_out_34734 = net_34734;
  assign seg_9_10_lutff_4_out_34736 = net_34736;
  assign seg_9_10_lutff_7_out_34739 = net_34739;
  assign seg_9_10_sp4_h_l_46_24008 = seg_8_10_sp4_h_r_46_24008;
  assign seg_9_10_sp4_h_r_12_34868 = net_34868;
  assign seg_9_10_sp4_h_r_2_38702 = net_38702;
  assign seg_9_10_sp4_r_v_b_41_38715 = net_38715;
  assign seg_9_11_lutff_5_out_34860 = net_34860;
  assign seg_9_11_sp4_h_r_10_38823 = net_38823;
  assign seg_9_12_sp4_h_r_34_31284 = seg_7_12_sp4_h_r_10_31284;
  assign seg_9_12_sp4_r_v_b_35_38843 = net_38843;
  assign seg_9_12_sp4_r_v_b_3_38589 = net_38589;
  assign seg_9_12_sp4_v_b_2_34759 = net_34759;
  assign seg_9_18_neigh_op_tnr_5_39675 = seg_10_19_lutff_5_out_39675;
  assign seg_9_18_neigh_op_tnr_6_39676 = seg_10_19_lutff_6_out_39676;
  assign seg_9_18_sp4_h_r_2_39686 = net_39686;
  assign seg_9_18_sp4_r_v_b_11_39335 = net_39335;
  assign seg_9_20_sp4_h_l_41_25241 = seg_5_20_sp4_h_r_4_25241;
  assign seg_9_20_sp4_v_b_6_35747 = seg_8_17_sp4_r_v_b_43_35747;
  assign seg_9_23_sp4_v_t_40_36605 = seg_8_25_sp4_r_v_b_29_36605;
  assign seg_9_27_lutff_1_out_36824 = net_36824;
  assign seg_9_27_lutff_5_out_36828 = net_36828;
  assign seg_9_27_lutff_7_out_36830 = net_36830;
  assign seg_9_27_neigh_op_rgt_2_40656 = seg_10_27_lutff_2_out_40656;
  assign seg_9_27_sp4_r_v_b_36_40801 = seg_10_29_sp4_v_b_12_40801;
  assign seg_9_28_lutff_2_out_36948 = net_36948;
  assign seg_9_28_lutff_5_out_36951 = net_36951;
  assign seg_9_28_neigh_op_bnr_7_40661 = seg_10_27_lutff_7_out_40661;
  assign seg_9_28_neigh_op_bot_5_36828 = seg_9_27_lutff_5_out_36828;
  assign seg_9_28_neigh_op_bot_7_36830 = seg_9_27_lutff_7_out_36830;
  assign seg_9_28_neigh_op_rgt_3_40780 = seg_10_28_lutff_3_out_40780;
  assign seg_9_28_neigh_op_top_5_37074 = seg_9_29_lutff_5_out_37074;
  assign seg_9_28_sp4_h_r_34_33252 = net_33252;
  assign seg_9_28_sp4_v_b_44_37101 = net_37101;
  assign seg_9_29_lutff_0_out_37069 = net_37069;
  assign seg_9_29_lutff_3_out_37072 = net_37072;
  assign seg_9_29_lutff_5_out_37074 = net_37074;
  assign seg_9_29_neigh_op_rgt_0_40900 = seg_10_29_lutff_0_out_40900;
  assign seg_9_29_neigh_op_rgt_5_40905 = seg_10_29_lutff_5_out_40905;
  assign seg_9_29_neigh_op_tnr_3_41026 = seg_10_30_lutff_3_out_41026;
  assign seg_9_29_neigh_op_tnr_4_41027 = seg_10_30_lutff_4_out_41027;
  assign seg_9_29_sp4_h_r_38_29568 = net_29568;
  assign seg_9_2_lutff_0_out_33712 = net_33712;
  assign seg_9_2_lutff_1_out_33713 = net_33713;
  assign seg_9_2_lutff_2_out_33714 = net_33714;
  assign seg_9_2_lutff_3_out_33715 = net_33715;
  assign seg_9_2_lutff_4_out_33716 = net_33716;
  assign seg_9_2_lutff_5_out_33717 = net_33717;
  assign seg_9_2_lutff_6_out_33718 = net_33718;
  assign seg_9_2_lutff_7_out_33719 = net_33719;
  assign seg_9_2_neigh_op_lft_3_29884 = seg_8_2_lutff_3_out_29884;
  assign seg_9_2_neigh_op_rgt_6_37549 = seg_10_2_lutff_6_out_37549;
  assign seg_9_2_neigh_op_rgt_7_37550 = seg_10_2_lutff_7_out_37550;
  assign seg_9_2_neigh_op_tnl_5_30045 = seg_8_3_lutff_5_out_30045;
  assign seg_9_2_neigh_op_tnr_2_37704 = seg_10_3_lutff_2_out_37704;
  assign seg_9_2_neigh_op_tnr_3_37705 = seg_10_3_lutff_3_out_37705;
  assign seg_9_2_neigh_op_tnr_4_37706 = seg_10_3_lutff_4_out_37706;
  assign seg_9_2_neigh_op_tnr_6_37708 = seg_10_3_lutff_6_out_37708;
  assign seg_9_2_neigh_op_top_1_33872 = seg_9_3_lutff_1_out_33872;
  assign seg_9_2_neigh_op_top_2_33873 = seg_9_3_lutff_2_out_33873;
  assign seg_9_2_neigh_op_top_4_33875 = seg_9_3_lutff_4_out_33875;
  assign seg_9_2_neigh_op_top_7_33878 = seg_9_3_lutff_7_out_33878;
  assign seg_9_2_sp4_v_b_27_33768 = seg_8_4_sp4_r_v_b_3_33768;
  assign seg_9_2_sp4_v_t_46_34028 = seg_8_4_sp4_r_v_b_35_34028;
  assign seg_9_30_lutff_0_out_37192 = net_37192;
  assign seg_9_30_lutff_5_out_37197 = net_37197;
  assign seg_9_30_lutff_7_out_37199 = net_37199;
  assign seg_9_30_neigh_op_bnr_0_40900 = seg_10_29_lutff_0_out_40900;
  assign seg_9_30_neigh_op_bnr_5_40905 = seg_10_29_lutff_5_out_40905;
  assign seg_9_30_neigh_op_rgt_3_41026 = seg_10_30_lutff_3_out_41026;
  assign seg_9_30_neigh_op_rgt_4_41027 = seg_10_30_lutff_4_out_41027;
  assign seg_9_30_neigh_op_tnl_6_33486 = seg_8_31_io_1_D_IN_0_33486;
  assign seg_9_30_sp4_v_b_20_37101 = seg_9_28_sp4_v_b_44_37101;
  assign seg_9_3_lutff_0_out_33871 = net_33871;
  assign seg_9_3_lutff_1_out_33872 = net_33872;
  assign seg_9_3_lutff_2_out_33873 = net_33873;
  assign seg_9_3_lutff_3_out_33874 = net_33874;
  assign seg_9_3_lutff_4_out_33875 = net_33875;
  assign seg_9_3_lutff_5_out_33876 = net_33876;
  assign seg_9_3_lutff_6_out_33877 = net_33877;
  assign seg_9_3_lutff_7_out_33878 = net_33878;
  assign seg_9_3_neigh_op_bnl_1_29882 = seg_8_2_lutff_1_out_29882;
  assign seg_9_3_neigh_op_bot_6_33718 = seg_9_2_lutff_6_out_33718;
  assign seg_9_3_neigh_op_lft_5_30045 = seg_8_3_lutff_5_out_30045;
  assign seg_9_3_neigh_op_top_5_33999 = seg_9_4_lutff_5_out_33999;
  assign seg_9_3_sp4_v_b_19_33774 = seg_8_3_sp4_r_v_b_19_33774;
  assign seg_9_4_lutff_1_out_33995 = net_33995;
  assign seg_9_4_lutff_5_out_33999 = net_33999;
  assign seg_9_4_neigh_op_bnl_5_30045 = seg_8_3_lutff_5_out_30045;
  assign seg_9_4_neigh_op_bot_0_33871 = seg_9_3_lutff_0_out_33871;
  assign seg_9_4_sp4_v_b_16_33899 = net_33899;
  assign seg_9_4_sp4_v_b_3_33768 = seg_8_4_sp4_r_v_b_3_33768;
  assign seg_9_5_neigh_op_bnl_1_30164 = seg_8_4_lutff_1_out_30164;
  assign seg_9_5_sp4_h_l_37_23390 = seg_5_5_sp4_h_r_0_23390;
  assign seg_9_5_sp4_r_v_b_23_37860 = net_37860;
  assign seg_9_5_sp4_v_b_5_33899 = seg_9_4_sp4_v_b_16_33899;
  assign seg_9_6_sp4_v_b_11_34028 = seg_8_4_sp4_r_v_b_35_34028;
  assign seg_9_8_lutff_5_out_34491 = net_34491;
  assign seg_9_8_lutff_6_out_34492 = net_34492;
  assign seg_9_8_lutff_7_out_34493 = net_34493;
  assign seg_9_8_neigh_op_rgt_2_38319 = seg_10_8_lutff_2_out_38319;
  assign seg_9_8_neigh_op_rgt_4_38321 = seg_10_8_lutff_4_out_38321;
  assign seg_9_8_neigh_op_rgt_6_38323 = seg_10_8_lutff_6_out_38323;
  assign seg_9_8_sp4_h_r_24_30790 = net_30790;
  assign seg_9_8_sp4_r_v_b_21_38227 = net_38227;
  assign seg_9_8_sp4_r_v_b_23_38229 = net_38229;
  assign seg_9_8_sp4_v_t_39_34759 = seg_9_12_sp4_v_b_2_34759;
  assign seg_9_9_sp4_h_r_10_38577 = seg_11_9_sp4_h_r_34_38577;
  wire gnd, vcc;
  GND gnd_cell (.Y(gnd));
  VCC vcc_cell (.Y(vcc));
  inout io_6_0_0;
  wire io_pad_6_0_0_din;
  wire io_pad_6_0_0_dout;
  wire io_pad_6_0_0_oe;
  IO_PAD io_pad_6_0_0 (
    .DIN(io_pad_6_0_0_din),
    .DOUT(io_pad_6_0_0_dout),
    .OE(io_pad_6_0_0_oe),
    .PACKAGEPIN(io_6_0_0)
  );
  inout io_7_0_0;
  wire io_pad_7_0_0_din;
  wire io_pad_7_0_0_dout;
  wire io_pad_7_0_0_oe;
  IO_PAD io_pad_7_0_0 (
    .DIN(io_pad_7_0_0_din),
    .DOUT(io_pad_7_0_0_dout),
    .OE(io_pad_7_0_0_oe),
    .PACKAGEPIN(io_7_0_0)
  );
  inout io_8_31_1;
  wire io_pad_8_31_1_din;
  wire io_pad_8_31_1_dout;
  wire io_pad_8_31_1_oe;
  IO_PAD io_pad_8_31_1 (
    .DIN(io_pad_8_31_1_din),
    .DOUT(io_pad_8_31_1_dout),
    .OE(io_pad_8_31_1_oe),
    .PACKAGEPIN(io_8_31_1)
  );
  inout io_12_31_1;
  wire io_pad_12_31_1_din;
  wire io_pad_12_31_1_dout;
  wire io_pad_12_31_1_oe;
  IO_PAD io_pad_12_31_1 (
    .DIN(io_pad_12_31_1_din),
    .DOUT(io_pad_12_31_1_dout),
    .OE(io_pad_12_31_1_oe),
    .PACKAGEPIN(io_12_31_1)
  );
  inout io_13_31_0;
  wire io_pad_13_31_0_din;
  wire io_pad_13_31_0_dout;
  wire io_pad_13_31_0_oe;
  IO_PAD io_pad_13_31_0 (
    .DIN(io_pad_13_31_0_din),
    .DOUT(io_pad_13_31_0_dout),
    .OE(io_pad_13_31_0_oe),
    .PACKAGEPIN(io_13_31_0)
  );
  inout io_17_0_0;
  wire io_pad_17_0_0_din;
  wire io_pad_17_0_0_dout;
  wire io_pad_17_0_0_oe;
  IO_PAD io_pad_17_0_0 (
    .DIN(io_pad_17_0_0_din),
    .DOUT(io_pad_17_0_0_dout),
    .OE(io_pad_17_0_0_oe),
    .PACKAGEPIN(io_17_0_0)
  );
  inout io_17_31_0;
  wire io_pad_17_31_0_din;
  wire io_pad_17_31_0_dout;
  wire io_pad_17_31_0_oe;
  IO_PAD io_pad_17_31_0 (
    .DIN(io_pad_17_31_0_din),
    .DOUT(io_pad_17_31_0_dout),
    .OE(io_pad_17_31_0_oe),
    .PACKAGEPIN(io_17_31_0)
  );
  inout io_18_0_0;
  wire io_pad_18_0_0_din;
  wire io_pad_18_0_0_dout;
  wire io_pad_18_0_0_oe;
  IO_PAD io_pad_18_0_0 (
    .DIN(io_pad_18_0_0_din),
    .DOUT(io_pad_18_0_0_dout),
    .OE(io_pad_18_0_0_oe),
    .PACKAGEPIN(io_18_0_0)
  );
  inout io_18_31_1;
  wire io_pad_18_31_1_din;
  wire io_pad_18_31_1_dout;
  wire io_pad_18_31_1_oe;
  IO_PAD io_pad_18_31_1 (
    .DIN(io_pad_18_31_1_din),
    .DOUT(io_pad_18_31_1_dout),
    .OE(io_pad_18_31_1_oe),
    .PACKAGEPIN(io_18_31_1)
  );
  inout io_22_0_1;
  wire io_pad_22_0_1_din;
  wire io_pad_22_0_1_dout;
  wire io_pad_22_0_1_oe;
  IO_PAD io_pad_22_0_1 (
    .DIN(io_pad_22_0_1_din),
    .DOUT(io_pad_22_0_1_dout),
    .OE(io_pad_22_0_1_oe),
    .PACKAGEPIN(io_22_0_1)
  );
  InMux inmux_10_10_42436_42481 (
    .I(net_42436),
    .O(net_42481)
  );
  InMux inmux_10_10_42441_42482 (
    .I(net_42441),
    .O(net_42482)
  );
  CEMux inmux_10_11_42560_42637 (
    .I(net_42560),
    .O(net_42637)
  );
  InMux inmux_10_11_42563_42618 (
    .I(net_42563),
    .O(net_42618)
  );
  InMux inmux_10_11_42576_42593 (
    .I(net_42576),
    .O(net_42593)
  );
  InMux inmux_10_11_42578_42605 (
    .I(net_42578),
    .O(net_42605)
  );
  InMux inmux_10_11_42581_42597 (
    .I(net_42581),
    .O(net_42597)
  );
  InMux inmux_10_11_42586_42606 (
    .I(net_42586),
    .O(net_42606)
  );
  InMux inmux_10_11_42587_42603 (
    .I(net_42587),
    .O(net_42603)
  );
  ClkMux inmux_10_11_5_42638 (
    .I(net_5),
    .O(net_42638)
  );
  InMux inmux_10_12_42681_42757 (
    .I(net_42681),
    .O(net_42757)
  );
  InMux inmux_10_12_42682_42727 (
    .I(net_42682),
    .O(net_42727)
  );
  InMux inmux_10_12_42684_42739 (
    .I(net_42684),
    .O(net_42739)
  );
  InMux inmux_10_12_42685_42740 (
    .I(net_42685),
    .O(net_42740)
  );
  InMux inmux_10_12_42686_42734 (
    .I(net_42686),
    .O(net_42734)
  );
  InMux inmux_10_12_42687_42745 (
    .I(net_42687),
    .O(net_42745)
  );
  InMux inmux_10_12_42689_42751 (
    .I(net_42689),
    .O(net_42751)
  );
  InMux inmux_10_12_42690_42716 (
    .I(net_42690),
    .O(net_42716)
  );
  InMux inmux_10_12_42692_42721 (
    .I(net_42692),
    .O(net_42721)
  );
  InMux inmux_10_12_42693_42715 (
    .I(net_42693),
    .O(net_42715)
  );
  InMux inmux_10_12_42696_42752 (
    .I(net_42696),
    .O(net_42752)
  );
  InMux inmux_10_12_42698_42758 (
    .I(net_42698),
    .O(net_42758)
  );
  CEMux inmux_10_12_42699_42760 (
    .I(net_42699),
    .O(net_42760)
  );
  InMux inmux_10_12_42700_42722 (
    .I(net_42700),
    .O(net_42722)
  );
  InMux inmux_10_12_42702_42746 (
    .I(net_42702),
    .O(net_42746)
  );
  InMux inmux_10_12_42703_42733 (
    .I(net_42703),
    .O(net_42733)
  );
  InMux inmux_10_12_42708_42728 (
    .I(net_42708),
    .O(net_42728)
  );
  InMux inmux_10_12_42713_42723 (
    .I(net_42713),
    .O(net_42723)
  );
  InMux inmux_10_12_42719_42729 (
    .I(net_42719),
    .O(net_42729)
  );
  InMux inmux_10_12_42725_42735 (
    .I(net_42725),
    .O(net_42735)
  );
  InMux inmux_10_12_42731_42741 (
    .I(net_42731),
    .O(net_42741)
  );
  InMux inmux_10_12_42737_42747 (
    .I(net_42737),
    .O(net_42747)
  );
  InMux inmux_10_12_42743_42753 (
    .I(net_42743),
    .O(net_42753)
  );
  InMux inmux_10_12_42749_42759 (
    .I(net_42749),
    .O(net_42759)
  );
  ClkMux inmux_10_12_5_42761 (
    .I(net_5),
    .O(net_42761)
  );
  InMux inmux_10_13_42799_42840 (
    .I(net_42799),
    .O(net_42840)
  );
  InMux inmux_10_13_42804_42851 (
    .I(net_42804),
    .O(net_42851)
  );
  InMux inmux_10_13_42805_42857 (
    .I(net_42805),
    .O(net_42857)
  );
  InMux inmux_10_13_42807_42838 (
    .I(net_42807),
    .O(net_42838)
  );
  InMux inmux_10_13_42808_42863 (
    .I(net_42808),
    .O(net_42863)
  );
  InMux inmux_10_13_42809_42845 (
    .I(net_42809),
    .O(net_42845)
  );
  InMux inmux_10_13_42810_42880 (
    .I(net_42810),
    .O(net_42880)
  );
  InMux inmux_10_13_42811_42874 (
    .I(net_42811),
    .O(net_42874)
  );
  InMux inmux_10_13_42812_42850 (
    .I(net_42812),
    .O(net_42850)
  );
  InMux inmux_10_13_42813_42868 (
    .I(net_42813),
    .O(net_42868)
  );
  InMux inmux_10_13_42815_42875 (
    .I(net_42815),
    .O(net_42875)
  );
  InMux inmux_10_13_42817_42856 (
    .I(net_42817),
    .O(net_42856)
  );
  InMux inmux_10_13_42822_42839 (
    .I(net_42822),
    .O(net_42839)
  );
  InMux inmux_10_13_42823_42869 (
    .I(net_42823),
    .O(net_42869)
  );
  InMux inmux_10_13_42828_42862 (
    .I(net_42828),
    .O(net_42862)
  );
  CEMux inmux_10_13_42831_42883 (
    .I(net_42831),
    .O(net_42883)
  );
  InMux inmux_10_13_42832_42881 (
    .I(net_42832),
    .O(net_42881)
  );
  InMux inmux_10_13_42835_42844 (
    .I(net_42835),
    .O(net_42844)
  );
  InMux inmux_10_13_42836_42846 (
    .I(net_42836),
    .O(net_42846)
  );
  InMux inmux_10_13_42842_42852 (
    .I(net_42842),
    .O(net_42852)
  );
  InMux inmux_10_13_42848_42858 (
    .I(net_42848),
    .O(net_42858)
  );
  InMux inmux_10_13_42854_42864 (
    .I(net_42854),
    .O(net_42864)
  );
  InMux inmux_10_13_42860_42870 (
    .I(net_42860),
    .O(net_42870)
  );
  InMux inmux_10_13_42866_42876 (
    .I(net_42866),
    .O(net_42876)
  );
  InMux inmux_10_13_42872_42882 (
    .I(net_42872),
    .O(net_42882)
  );
  ClkMux inmux_10_13_5_42884 (
    .I(net_5),
    .O(net_42884)
  );
  InMux inmux_10_14_42927_43003 (
    .I(net_42927),
    .O(net_43003)
  );
  InMux inmux_10_14_42936_42984 (
    .I(net_42936),
    .O(net_42984)
  );
  InMux inmux_10_14_42938_42998 (
    .I(net_42938),
    .O(net_42998)
  );
  InMux inmux_10_14_42941_42992 (
    .I(net_42941),
    .O(net_42992)
  );
  InMux inmux_10_14_42942_42974 (
    .I(net_42942),
    .O(net_42974)
  );
  InMux inmux_10_14_42945_42962 (
    .I(net_42945),
    .O(net_42962)
  );
  InMux inmux_10_14_42947_42969 (
    .I(net_42947),
    .O(net_42969)
  );
  InMux inmux_10_14_42958_42981 (
    .I(net_42958),
    .O(net_42981)
  );
  ClkMux inmux_10_14_5_43007 (
    .I(net_5),
    .O(net_43007)
  );
  CEMux inmux_10_14_6_43006 (
    .I(net_6),
    .O(net_43006)
  );
  InMux inmux_10_15_43052_43109 (
    .I(net_43052),
    .O(net_43109)
  );
  InMux inmux_10_15_43056_43085 (
    .I(net_43056),
    .O(net_43085)
  );
  InMux inmux_10_15_43074_43096 (
    .I(net_43074),
    .O(net_43096)
  );
  ClkMux inmux_10_15_5_43130 (
    .I(net_5),
    .O(net_43130)
  );
  CEMux inmux_10_15_6_43129 (
    .I(net_6),
    .O(net_43129)
  );
  InMux inmux_10_17_43300_43355 (
    .I(net_43300),
    .O(net_43355)
  );
  InMux inmux_10_17_43302_43367 (
    .I(net_43302),
    .O(net_43367)
  );
  InMux inmux_10_17_43309_43336 (
    .I(net_43309),
    .O(net_43336)
  );
  InMux inmux_10_17_43311_43372 (
    .I(net_43311),
    .O(net_43372)
  );
  InMux inmux_10_17_43315_43349 (
    .I(net_43315),
    .O(net_43349)
  );
  InMux inmux_10_17_43321_43331 (
    .I(net_43321),
    .O(net_43331)
  );
  InMux inmux_10_17_43322_43342 (
    .I(net_43322),
    .O(net_43342)
  );
  InMux inmux_10_17_43325_43360 (
    .I(net_43325),
    .O(net_43360)
  );
  InMux inmux_10_17_43334_43344 (
    .I(net_43334),
    .O(net_43344)
  );
  InMux inmux_10_17_43340_43350 (
    .I(net_43340),
    .O(net_43350)
  );
  InMux inmux_10_17_43346_43356 (
    .I(net_43346),
    .O(net_43356)
  );
  InMux inmux_10_17_43352_43362 (
    .I(net_43352),
    .O(net_43362)
  );
  InMux inmux_10_17_43358_43368 (
    .I(net_43358),
    .O(net_43368)
  );
  InMux inmux_10_17_43364_43374 (
    .I(net_43364),
    .O(net_43374)
  );
  ClkMux inmux_10_17_5_43376 (
    .I(net_5),
    .O(net_43376)
  );
  InMux inmux_10_18_43414_43455 (
    .I(net_43414),
    .O(net_43455)
  );
  InMux inmux_10_18_43424_43484 (
    .I(net_43424),
    .O(net_43484)
  );
  InMux inmux_10_18_43430_43471 (
    .I(net_43430),
    .O(net_43471)
  );
  InMux inmux_10_18_43436_43460 (
    .I(net_43436),
    .O(net_43460)
  );
  InMux inmux_10_18_43437_43466 (
    .I(net_43437),
    .O(net_43466)
  );
  InMux inmux_10_18_43441_43490 (
    .I(net_43441),
    .O(net_43490)
  );
  InMux inmux_10_18_43443_43453 (
    .I(net_43443),
    .O(net_43453)
  );
  InMux inmux_10_18_43447_43477 (
    .I(net_43447),
    .O(net_43477)
  );
  InMux inmux_10_18_43450_43495 (
    .I(net_43450),
    .O(net_43495)
  );
  InMux inmux_10_18_43451_43461 (
    .I(net_43451),
    .O(net_43461)
  );
  InMux inmux_10_18_43457_43467 (
    .I(net_43457),
    .O(net_43467)
  );
  InMux inmux_10_18_43463_43473 (
    .I(net_43463),
    .O(net_43473)
  );
  InMux inmux_10_18_43469_43479 (
    .I(net_43469),
    .O(net_43479)
  );
  InMux inmux_10_18_43475_43485 (
    .I(net_43475),
    .O(net_43485)
  );
  InMux inmux_10_18_43481_43491 (
    .I(net_43481),
    .O(net_43491)
  );
  InMux inmux_10_18_43487_43497 (
    .I(net_43487),
    .O(net_43497)
  );
  ClkMux inmux_10_18_5_43499 (
    .I(net_5),
    .O(net_43499)
  );
  InMux inmux_10_19_43537_43578 (
    .I(net_43537),
    .O(net_43578)
  );
  InMux inmux_10_19_43544_43589 (
    .I(net_43544),
    .O(net_43589)
  );
  InMux inmux_10_19_43548_43613 (
    .I(net_43548),
    .O(net_43613)
  );
  InMux inmux_10_19_43549_43619 (
    .I(net_43549),
    .O(net_43619)
  );
  InMux inmux_10_19_43550_43576 (
    .I(net_43550),
    .O(net_43576)
  );
  InMux inmux_10_19_43551_43582 (
    .I(net_43551),
    .O(net_43582)
  );
  InMux inmux_10_19_43554_43600 (
    .I(net_43554),
    .O(net_43600)
  );
  InMux inmux_10_19_43569_43594 (
    .I(net_43569),
    .O(net_43594)
  );
  InMux inmux_10_19_43571_43606 (
    .I(net_43571),
    .O(net_43606)
  );
  InMux inmux_10_19_43574_43584 (
    .I(net_43574),
    .O(net_43584)
  );
  InMux inmux_10_19_43580_43590 (
    .I(net_43580),
    .O(net_43590)
  );
  InMux inmux_10_19_43586_43596 (
    .I(net_43586),
    .O(net_43596)
  );
  InMux inmux_10_19_43592_43602 (
    .I(net_43592),
    .O(net_43602)
  );
  InMux inmux_10_19_43598_43608 (
    .I(net_43598),
    .O(net_43608)
  );
  InMux inmux_10_19_43604_43614 (
    .I(net_43604),
    .O(net_43614)
  );
  InMux inmux_10_19_43610_43620 (
    .I(net_43610),
    .O(net_43620)
  );
  ClkMux inmux_10_19_5_43622 (
    .I(net_5),
    .O(net_43622)
  );
  InMux inmux_10_20_43660_43701 (
    .I(net_43660),
    .O(net_43701)
  );
  InMux inmux_10_20_43666_43706 (
    .I(net_43666),
    .O(net_43706)
  );
  InMux inmux_10_20_43668_43718 (
    .I(net_43668),
    .O(net_43718)
  );
  InMux inmux_10_20_43673_43699 (
    .I(net_43673),
    .O(net_43699)
  );
  InMux inmux_10_20_43691_43711 (
    .I(net_43691),
    .O(net_43711)
  );
  InMux inmux_10_20_43697_43707 (
    .I(net_43697),
    .O(net_43707)
  );
  InMux inmux_10_20_43703_43713 (
    .I(net_43703),
    .O(net_43713)
  );
  InMux inmux_10_20_43709_43719 (
    .I(net_43709),
    .O(net_43719)
  );
  ClkMux inmux_10_20_5_43745 (
    .I(net_5),
    .O(net_43745)
  );
  InMux inmux_10_26_44413_44451 (
    .I(net_44413),
    .O(net_44451)
  );
  InMux inmux_10_26_44413_44478 (
    .I(net_44413),
    .O(net_44478)
  );
  CEMux inmux_10_26_44430_44482 (
    .I(net_44430),
    .O(net_44482)
  );
  InMux inmux_10_26_44434_44448 (
    .I(net_44434),
    .O(net_44448)
  );
  ClkMux inmux_10_26_5_44483 (
    .I(net_5),
    .O(net_44483)
  );
  InMux inmux_10_27_44529_44567 (
    .I(net_44529),
    .O(net_44567)
  );
  InMux inmux_10_27_44531_44572 (
    .I(net_44531),
    .O(net_44572)
  );
  InMux inmux_10_27_44532_44590 (
    .I(net_44532),
    .O(net_44590)
  );
  InMux inmux_10_27_44533_44584 (
    .I(net_44533),
    .O(net_44584)
  );
  InMux inmux_10_27_44537_44604 (
    .I(net_44537),
    .O(net_44604)
  );
  InMux inmux_10_27_44539_44595 (
    .I(net_44539),
    .O(net_44595)
  );
  InMux inmux_10_27_44541_44561 (
    .I(net_44541),
    .O(net_44561)
  );
  InMux inmux_10_27_44549_44579 (
    .I(net_44549),
    .O(net_44579)
  );
  CEMux inmux_10_27_44553_44605 (
    .I(net_44553),
    .O(net_44605)
  );
  InMux inmux_10_27_44554_44596 (
    .I(net_44554),
    .O(net_44596)
  );
  InMux inmux_10_27_44554_44601 (
    .I(net_44554),
    .O(net_44601)
  );
  InMux inmux_10_27_44564_44574 (
    .I(net_44564),
    .O(net_44574)
  );
  InMux inmux_10_27_44570_44580 (
    .I(net_44570),
    .O(net_44580)
  );
  InMux inmux_10_27_44576_44586 (
    .I(net_44576),
    .O(net_44586)
  );
  InMux inmux_10_27_44582_44592 (
    .I(net_44582),
    .O(net_44592)
  );
  ClkMux inmux_10_27_5_44606 (
    .I(net_5),
    .O(net_44606)
  );
  InMux inmux_10_28_44653_44727 (
    .I(net_44653),
    .O(net_44727)
  );
  InMux inmux_10_28_44655_44694 (
    .I(net_44655),
    .O(net_44694)
  );
  InMux inmux_10_28_44656_44697 (
    .I(net_44656),
    .O(net_44697)
  );
  InMux inmux_10_28_44660_44701 (
    .I(net_44660),
    .O(net_44701)
  );
  InMux inmux_10_28_44660_44713 (
    .I(net_44660),
    .O(net_44713)
  );
  InMux inmux_10_28_44663_44702 (
    .I(net_44663),
    .O(net_44702)
  );
  InMux inmux_10_28_44663_44712 (
    .I(net_44663),
    .O(net_44712)
  );
  InMux inmux_10_28_44663_44726 (
    .I(net_44663),
    .O(net_44726)
  );
  InMux inmux_10_28_44664_44696 (
    .I(net_44664),
    .O(net_44696)
  );
  InMux inmux_10_28_44670_44695 (
    .I(net_44670),
    .O(net_44695)
  );
  InMux inmux_10_28_44675_44714 (
    .I(net_44675),
    .O(net_44714)
  );
  CEMux inmux_10_28_44676_44728 (
    .I(net_44676),
    .O(net_44728)
  );
  InMux inmux_10_28_44680_44703 (
    .I(net_44680),
    .O(net_44703)
  );
  InMux inmux_10_28_44680_44715 (
    .I(net_44680),
    .O(net_44715)
  );
  ClkMux inmux_10_28_5_44729 (
    .I(net_5),
    .O(net_44729)
  );
  InMux inmux_10_29_44773_44818 (
    .I(net_44773),
    .O(net_44818)
  );
  InMux inmux_10_29_44773_44825 (
    .I(net_44773),
    .O(net_44825)
  );
  CEMux inmux_10_29_44774_44851 (
    .I(net_44774),
    .O(net_44851)
  );
  InMux inmux_10_29_44783_44807 (
    .I(net_44783),
    .O(net_44807)
  );
  InMux inmux_10_29_44783_44824 (
    .I(net_44783),
    .O(net_44824)
  );
  InMux inmux_10_29_44783_44836 (
    .I(net_44783),
    .O(net_44836)
  );
  InMux inmux_10_29_44783_44841 (
    .I(net_44783),
    .O(net_44841)
  );
  InMux inmux_10_29_44783_44848 (
    .I(net_44783),
    .O(net_44848)
  );
  InMux inmux_10_29_44784_44806 (
    .I(net_44784),
    .O(net_44806)
  );
  InMux inmux_10_29_44784_44823 (
    .I(net_44784),
    .O(net_44823)
  );
  InMux inmux_10_29_44784_44835 (
    .I(net_44784),
    .O(net_44835)
  );
  InMux inmux_10_29_44784_44844 (
    .I(net_44784),
    .O(net_44844)
  );
  InMux inmux_10_29_44784_44847 (
    .I(net_44784),
    .O(net_44847)
  );
  InMux inmux_10_29_44788_44805 (
    .I(net_44788),
    .O(net_44805)
  );
  InMux inmux_10_29_44788_44826 (
    .I(net_44788),
    .O(net_44826)
  );
  InMux inmux_10_29_44788_44838 (
    .I(net_44788),
    .O(net_44838)
  );
  InMux inmux_10_29_44788_44843 (
    .I(net_44788),
    .O(net_44843)
  );
  InMux inmux_10_29_44788_44850 (
    .I(net_44788),
    .O(net_44850)
  );
  InMux inmux_10_29_44793_44808 (
    .I(net_44793),
    .O(net_44808)
  );
  InMux inmux_10_29_44793_44837 (
    .I(net_44793),
    .O(net_44837)
  );
  InMux inmux_10_29_44793_44842 (
    .I(net_44793),
    .O(net_44842)
  );
  InMux inmux_10_29_44793_44849 (
    .I(net_44793),
    .O(net_44849)
  );
  InMux inmux_10_29_44803_44817 (
    .I(net_44803),
    .O(net_44817)
  );
  ClkMux inmux_10_29_5_44852 (
    .I(net_5),
    .O(net_44852)
  );
  InMux inmux_10_2_41453_41515 (
    .I(net_41453),
    .O(net_41515)
  );
  InMux inmux_10_2_41454_41485 (
    .I(net_41454),
    .O(net_41485)
  );
  InMux inmux_10_2_41455_41520 (
    .I(net_41455),
    .O(net_41520)
  );
  InMux inmux_10_2_41455_41529 (
    .I(net_41455),
    .O(net_41529)
  );
  InMux inmux_10_2_41457_41491 (
    .I(net_41457),
    .O(net_41491)
  );
  InMux inmux_10_2_41458_41497 (
    .I(net_41458),
    .O(net_41497)
  );
  CEMux inmux_10_2_41462_41530 (
    .I(net_41462),
    .O(net_41530)
  );
  InMux inmux_10_2_41463_41504 (
    .I(net_41463),
    .O(net_41504)
  );
  InMux inmux_10_2_41465_41509 (
    .I(net_41465),
    .O(net_41509)
  );
  InMux inmux_10_2_41471_41522 (
    .I(net_41471),
    .O(net_41522)
  );
  InMux inmux_10_2_41477_41526 (
    .I(net_41477),
    .O(net_41526)
  );
  InMux inmux_10_2_41489_41499 (
    .I(net_41489),
    .O(net_41499)
  );
  InMux inmux_10_2_41495_41505 (
    .I(net_41495),
    .O(net_41505)
  );
  InMux inmux_10_2_41501_41511 (
    .I(net_41501),
    .O(net_41511)
  );
  InMux inmux_10_2_41507_41517 (
    .I(net_41507),
    .O(net_41517)
  );
  ClkMux inmux_10_2_5_41531 (
    .I(net_5),
    .O(net_41531)
  );
  InMux inmux_10_30_44895_44930 (
    .I(net_44895),
    .O(net_44930)
  );
  CEMux inmux_10_30_44897_44974 (
    .I(net_44897),
    .O(net_44974)
  );
  InMux inmux_10_30_44899_44966 (
    .I(net_44899),
    .O(net_44966)
  );
  InMux inmux_10_30_44900_44929 (
    .I(net_44900),
    .O(net_44929)
  );
  InMux inmux_10_30_44900_44965 (
    .I(net_44900),
    .O(net_44965)
  );
  InMux inmux_10_30_44903_44941 (
    .I(net_44903),
    .O(net_44941)
  );
  InMux inmux_10_30_44903_44972 (
    .I(net_44903),
    .O(net_44972)
  );
  InMux inmux_10_30_44905_44946 (
    .I(net_44905),
    .O(net_44946)
  );
  InMux inmux_10_30_44905_44953 (
    .I(net_44905),
    .O(net_44953)
  );
  InMux inmux_10_30_44907_44943 (
    .I(net_44907),
    .O(net_44943)
  );
  InMux inmux_10_30_44907_44948 (
    .I(net_44907),
    .O(net_44948)
  );
  InMux inmux_10_30_44907_44955 (
    .I(net_44907),
    .O(net_44955)
  );
  InMux inmux_10_30_44908_44940 (
    .I(net_44908),
    .O(net_44940)
  );
  InMux inmux_10_30_44908_44971 (
    .I(net_44908),
    .O(net_44971)
  );
  InMux inmux_10_30_44911_44942 (
    .I(net_44911),
    .O(net_44942)
  );
  InMux inmux_10_30_44913_44949 (
    .I(net_44913),
    .O(net_44949)
  );
  InMux inmux_10_30_44917_44952 (
    .I(net_44917),
    .O(net_44952)
  );
  InMux inmux_10_30_44917_44973 (
    .I(net_44917),
    .O(net_44973)
  );
  InMux inmux_10_30_44922_44947 (
    .I(net_44922),
    .O(net_44947)
  );
  InMux inmux_10_30_44922_44964 (
    .I(net_44922),
    .O(net_44964)
  );
  InMux inmux_10_30_44923_44970 (
    .I(net_44923),
    .O(net_44970)
  );
  InMux inmux_10_30_44925_44967 (
    .I(net_44925),
    .O(net_44967)
  );
  InMux inmux_10_30_44926_44954 (
    .I(net_44926),
    .O(net_44954)
  );
  ClkMux inmux_10_30_5_44975 (
    .I(net_5),
    .O(net_44975)
  );
  CEMux inmux_10_3_41576_41653 (
    .I(net_41576),
    .O(net_41653)
  );
  InMux inmux_10_3_41585_41633 (
    .I(net_41585),
    .O(net_41633)
  );
  InMux inmux_10_3_41587_41619 (
    .I(net_41587),
    .O(net_41619)
  );
  InMux inmux_10_3_41588_41644 (
    .I(net_41588),
    .O(net_41644)
  );
  InMux inmux_10_3_41594_41621 (
    .I(net_41594),
    .O(net_41621)
  );
  InMux inmux_10_3_41594_41628 (
    .I(net_41594),
    .O(net_41628)
  );
  InMux inmux_10_3_41594_41631 (
    .I(net_41594),
    .O(net_41631)
  );
  InMux inmux_10_3_41594_41643 (
    .I(net_41594),
    .O(net_41643)
  );
  InMux inmux_10_3_41600_41651 (
    .I(net_41600),
    .O(net_41651)
  );
  InMux inmux_10_3_41601_41645 (
    .I(net_41601),
    .O(net_41645)
  );
  InMux inmux_10_3_41601_41652 (
    .I(net_41601),
    .O(net_41652)
  );
  InMux inmux_10_3_41605_41626 (
    .I(net_41605),
    .O(net_41626)
  );
  ClkMux inmux_10_3_5_41654 (
    .I(net_5),
    .O(net_41654)
  );
  InMux inmux_10_7_42071_42129 (
    .I(net_42071),
    .O(net_42129)
  );
  InMux inmux_10_7_42082_42132 (
    .I(net_42082),
    .O(net_42132)
  );
  InMux inmux_10_8_42192_42242 (
    .I(net_42192),
    .O(net_42242)
  );
  InMux inmux_10_8_42192_42264 (
    .I(net_42192),
    .O(net_42264)
  );
  InMux inmux_10_8_42194_42223 (
    .I(net_42194),
    .O(net_42223)
  );
  InMux inmux_10_8_42195_42224 (
    .I(net_42195),
    .O(net_42224)
  );
  InMux inmux_10_8_42196_42240 (
    .I(net_42196),
    .O(net_42240)
  );
  InMux inmux_10_8_42197_42230 (
    .I(net_42197),
    .O(net_42230)
  );
  InMux inmux_10_8_42200_42231 (
    .I(net_42200),
    .O(net_42231)
  );
  InMux inmux_10_8_42200_42258 (
    .I(net_42200),
    .O(net_42258)
  );
  InMux inmux_10_8_42203_42266 (
    .I(net_42203),
    .O(net_42266)
  );
  InMux inmux_10_8_42205_42229 (
    .I(net_42205),
    .O(net_42229)
  );
  InMux inmux_10_8_42205_42246 (
    .I(net_42205),
    .O(net_42246)
  );
  InMux inmux_10_8_42209_42222 (
    .I(net_42209),
    .O(net_42222)
  );
  InMux inmux_10_8_42209_42243 (
    .I(net_42209),
    .O(net_42243)
  );
  InMux inmux_10_8_42209_42267 (
    .I(net_42209),
    .O(net_42267)
  );
  InMux inmux_10_8_42210_42225 (
    .I(net_42210),
    .O(net_42225)
  );
  InMux inmux_10_8_42211_42265 (
    .I(net_42211),
    .O(net_42265)
  );
  InMux inmux_10_8_42212_42228 (
    .I(net_42212),
    .O(net_42228)
  );
  InMux inmux_10_8_42212_42237 (
    .I(net_42212),
    .O(net_42237)
  );
  CEMux inmux_10_8_42216_42268 (
    .I(net_42216),
    .O(net_42268)
  );
  InMux inmux_10_8_42220_42241 (
    .I(net_42220),
    .O(net_42241)
  );
  ClkMux inmux_10_8_5_42269 (
    .I(net_5),
    .O(net_42269)
  );
  CEMux inmux_11_10_46268_46345 (
    .I(net_46268),
    .O(net_46345)
  );
  InMux inmux_11_10_46269_46338 (
    .I(net_46269),
    .O(net_46338)
  );
  InMux inmux_11_10_46271_46300 (
    .I(net_46271),
    .O(net_46300)
  );
  InMux inmux_11_10_46271_46319 (
    .I(net_46271),
    .O(net_46319)
  );
  InMux inmux_11_10_46273_46336 (
    .I(net_46273),
    .O(net_46336)
  );
  InMux inmux_11_10_46273_46341 (
    .I(net_46273),
    .O(net_46341)
  );
  InMux inmux_11_10_46276_46302 (
    .I(net_46276),
    .O(net_46302)
  );
  InMux inmux_11_10_46277_46337 (
    .I(net_46277),
    .O(net_46337)
  );
  InMux inmux_11_10_46277_46342 (
    .I(net_46277),
    .O(net_46342)
  );
  InMux inmux_11_10_46279_46301 (
    .I(net_46279),
    .O(net_46301)
  );
  SRMux inmux_11_10_46286_46347 (
    .I(net_46286),
    .O(net_46347)
  );
  InMux inmux_11_10_46292_46324 (
    .I(net_46292),
    .O(net_46324)
  );
  InMux inmux_11_10_46292_46331 (
    .I(net_46292),
    .O(net_46331)
  );
  InMux inmux_11_10_46294_46317 (
    .I(net_46294),
    .O(net_46317)
  );
  InMux inmux_11_10_46294_46329 (
    .I(net_46294),
    .O(net_46329)
  );
  InMux inmux_11_10_46297_46299 (
    .I(net_46297),
    .O(net_46299)
  );
  ClkMux inmux_11_10_5_46346 (
    .I(net_5),
    .O(net_46346)
  );
  InMux inmux_11_11_46407_46436 (
    .I(net_46407),
    .O(net_46436)
  );
  InMux inmux_11_11_46419_46464 (
    .I(net_46419),
    .O(net_46464)
  );
  ClkMux inmux_11_11_5_46469 (
    .I(net_5),
    .O(net_46469)
  );
  CEMux inmux_11_11_6_46468 (
    .I(net_6),
    .O(net_46468)
  );
  InMux inmux_11_12_46513_46563 (
    .I(net_46513),
    .O(net_46563)
  );
  InMux inmux_11_12_46514_46581 (
    .I(net_46514),
    .O(net_46581)
  );
  InMux inmux_11_12_46517_46572 (
    .I(net_46517),
    .O(net_46572)
  );
  InMux inmux_11_12_46519_46551 (
    .I(net_46519),
    .O(net_46551)
  );
  InMux inmux_11_12_46525_46557 (
    .I(net_46525),
    .O(net_46557)
  );
  InMux inmux_11_12_46529_46565 (
    .I(net_46529),
    .O(net_46565)
  );
  InMux inmux_11_12_46532_46588 (
    .I(net_46532),
    .O(net_46588)
  );
  InMux inmux_11_12_46533_46570 (
    .I(net_46533),
    .O(net_46570)
  );
  InMux inmux_11_12_46534_46552 (
    .I(net_46534),
    .O(net_46552)
  );
  InMux inmux_11_12_46534_46566 (
    .I(net_46534),
    .O(net_46566)
  );
  InMux inmux_11_12_46534_46571 (
    .I(net_46534),
    .O(net_46571)
  );
  InMux inmux_11_12_46535_46553 (
    .I(net_46535),
    .O(net_46553)
  );
  InMux inmux_11_12_46537_46554 (
    .I(net_46537),
    .O(net_46554)
  );
  InMux inmux_11_12_46537_46564 (
    .I(net_46537),
    .O(net_46564)
  );
  InMux inmux_11_12_46537_46569 (
    .I(net_46537),
    .O(net_46569)
  );
  ClkMux inmux_11_12_5_46592 (
    .I(net_5),
    .O(net_46592)
  );
  CEMux inmux_11_12_6_46591 (
    .I(net_6),
    .O(net_46591)
  );
  InMux inmux_11_13_46639_46704 (
    .I(net_46639),
    .O(net_46704)
  );
  InMux inmux_11_13_46640_46669 (
    .I(net_46640),
    .O(net_46669)
  );
  InMux inmux_11_13_46640_46676 (
    .I(net_46640),
    .O(net_46676)
  );
  InMux inmux_11_13_46640_46681 (
    .I(net_46640),
    .O(net_46681)
  );
  InMux inmux_11_13_46640_46693 (
    .I(net_46640),
    .O(net_46693)
  );
  InMux inmux_11_13_46640_46698 (
    .I(net_46640),
    .O(net_46698)
  );
  InMux inmux_11_13_46640_46707 (
    .I(net_46640),
    .O(net_46707)
  );
  InMux inmux_11_13_46641_46701 (
    .I(net_46641),
    .O(net_46701)
  );
  InMux inmux_11_13_46642_46712 (
    .I(net_46642),
    .O(net_46712)
  );
  InMux inmux_11_13_46644_46682 (
    .I(net_46644),
    .O(net_46682)
  );
  InMux inmux_11_13_46645_46671 (
    .I(net_46645),
    .O(net_46671)
  );
  InMux inmux_11_13_46646_46670 (
    .I(net_46646),
    .O(net_46670)
  );
  InMux inmux_11_13_46646_46675 (
    .I(net_46646),
    .O(net_46675)
  );
  InMux inmux_11_13_46646_46680 (
    .I(net_46646),
    .O(net_46680)
  );
  InMux inmux_11_13_46646_46694 (
    .I(net_46646),
    .O(net_46694)
  );
  InMux inmux_11_13_46646_46699 (
    .I(net_46646),
    .O(net_46699)
  );
  InMux inmux_11_13_46646_46706 (
    .I(net_46646),
    .O(net_46706)
  );
  InMux inmux_11_13_46647_46688 (
    .I(net_46647),
    .O(net_46688)
  );
  InMux inmux_11_13_46648_46692 (
    .I(net_46648),
    .O(net_46692)
  );
  InMux inmux_11_13_46650_46677 (
    .I(net_46650),
    .O(net_46677)
  );
  InMux inmux_11_13_46652_46683 (
    .I(net_46652),
    .O(net_46683)
  );
  InMux inmux_11_13_46653_46668 (
    .I(net_46653),
    .O(net_46668)
  );
  InMux inmux_11_13_46656_46695 (
    .I(net_46656),
    .O(net_46695)
  );
  InMux inmux_11_13_46658_46674 (
    .I(net_46658),
    .O(net_46674)
  );
  InMux inmux_11_13_46663_46705 (
    .I(net_46663),
    .O(net_46705)
  );
  InMux inmux_11_13_46665_46700 (
    .I(net_46665),
    .O(net_46700)
  );
  InMux inmux_11_14_46758_46815 (
    .I(net_46758),
    .O(net_46815)
  );
  InMux inmux_11_14_46760_46829 (
    .I(net_46760),
    .O(net_46829)
  );
  InMux inmux_11_14_46762_46836 (
    .I(net_46762),
    .O(net_46836)
  );
  InMux inmux_11_14_46764_46798 (
    .I(net_46764),
    .O(net_46798)
  );
  InMux inmux_11_14_46765_46794 (
    .I(net_46765),
    .O(net_46794)
  );
  InMux inmux_11_14_46768_46821 (
    .I(net_46768),
    .O(net_46821)
  );
  InMux inmux_11_14_46768_46833 (
    .I(net_46768),
    .O(net_46833)
  );
  InMux inmux_11_14_46769_46800 (
    .I(net_46769),
    .O(net_46800)
  );
  InMux inmux_11_14_46773_46822 (
    .I(net_46773),
    .O(net_46822)
  );
  InMux inmux_11_14_46774_46805 (
    .I(net_46774),
    .O(net_46805)
  );
  InMux inmux_11_14_46774_46824 (
    .I(net_46774),
    .O(net_46824)
  );
  CEMux inmux_11_14_46776_46837 (
    .I(net_46776),
    .O(net_46837)
  );
  InMux inmux_11_14_46780_46812 (
    .I(net_46780),
    .O(net_46812)
  );
  InMux inmux_11_14_46780_46834 (
    .I(net_46780),
    .O(net_46834)
  );
  InMux inmux_11_14_46784_46823 (
    .I(net_46784),
    .O(net_46823)
  );
  InMux inmux_11_14_46784_46835 (
    .I(net_46784),
    .O(net_46835)
  );
  ClkMux inmux_11_14_5_46838 (
    .I(net_5),
    .O(net_46838)
  );
  InMux inmux_11_15_46884_46951 (
    .I(net_46884),
    .O(net_46951)
  );
  CEMux inmux_11_15_46892_46960 (
    .I(net_46892),
    .O(net_46960)
  );
  InMux inmux_11_15_46894_46940 (
    .I(net_46894),
    .O(net_46940)
  );
  InMux inmux_11_15_46898_46927 (
    .I(net_46898),
    .O(net_46927)
  );
  InMux inmux_11_15_46905_46932 (
    .I(net_46905),
    .O(net_46932)
  );
  ClkMux inmux_11_15_5_46961 (
    .I(net_5),
    .O(net_46961)
  );
  CEMux inmux_11_16_47006_47083 (
    .I(net_47006),
    .O(net_47083)
  );
  InMux inmux_11_16_47009_47069 (
    .I(net_47009),
    .O(net_47069)
  );
  ClkMux inmux_11_16_5_47084 (
    .I(net_5),
    .O(net_47084)
  );
  InMux inmux_11_17_47128_47166 (
    .I(net_47128),
    .O(net_47166)
  );
  InMux inmux_11_17_47148_47168 (
    .I(net_47148),
    .O(net_47168)
  );
  ClkMux inmux_11_17_5_47207 (
    .I(net_5),
    .O(net_47207)
  );
  InMux inmux_11_18_47252_47290 (
    .I(net_47252),
    .O(net_47290)
  );
  InMux inmux_11_18_47252_47297 (
    .I(net_47252),
    .O(net_47297)
  );
  InMux inmux_11_18_47258_47289 (
    .I(net_47258),
    .O(net_47289)
  );
  CEMux inmux_11_18_47268_47329 (
    .I(net_47268),
    .O(net_47329)
  );
  InMux inmux_11_18_47269_47291 (
    .I(net_47269),
    .O(net_47291)
  );
  InMux inmux_11_18_47271_47298 (
    .I(net_47271),
    .O(net_47298)
  );
  InMux inmux_11_18_47272_47304 (
    .I(net_47272),
    .O(net_47304)
  );
  InMux inmux_11_18_47274_47308 (
    .I(net_47274),
    .O(net_47308)
  );
  InMux inmux_11_18_47275_47292 (
    .I(net_47275),
    .O(net_47292)
  );
  InMux inmux_11_18_47275_47295 (
    .I(net_47275),
    .O(net_47295)
  );
  InMux inmux_11_18_47276_47296 (
    .I(net_47276),
    .O(net_47296)
  );
  InMux inmux_11_18_47279_47314 (
    .I(net_47279),
    .O(net_47314)
  );
  ClkMux inmux_11_18_5_47330 (
    .I(net_5),
    .O(net_47330)
  );
  InMux inmux_11_19_47374_47424 (
    .I(net_47374),
    .O(net_47424)
  );
  InMux inmux_11_19_47377_47418 (
    .I(net_47377),
    .O(net_47418)
  );
  InMux inmux_11_19_47382_47420 (
    .I(net_47382),
    .O(net_47420)
  );
  InMux inmux_11_19_47385_47445 (
    .I(net_47385),
    .O(net_47445)
  );
  CEMux inmux_11_19_47391_47452 (
    .I(net_47391),
    .O(net_47452)
  );
  InMux inmux_11_19_47397_47419 (
    .I(net_47397),
    .O(net_47419)
  );
  InMux inmux_11_19_47403_47421 (
    .I(net_47403),
    .O(net_47421)
  );
  ClkMux inmux_11_19_5_47453 (
    .I(net_5),
    .O(net_47453)
  );
  InMux inmux_11_20_47498_47543 (
    .I(net_47498),
    .O(net_47543)
  );
  InMux inmux_11_20_47505_47565 (
    .I(net_47505),
    .O(net_47565)
  );
  InMux inmux_11_20_47516_47538 (
    .I(net_47516),
    .O(net_47538)
  );
  ClkMux inmux_11_20_5_47576 (
    .I(net_5),
    .O(net_47576)
  );
  CEMux inmux_11_20_6_47575 (
    .I(net_6),
    .O(net_47575)
  );
  CEMux inmux_11_23_47883_47944 (
    .I(net_47883),
    .O(net_47944)
  );
  InMux inmux_11_23_47892_47936 (
    .I(net_47892),
    .O(net_47936)
  );
  ClkMux inmux_11_23_5_47945 (
    .I(net_5),
    .O(net_47945)
  );
  InMux inmux_11_29_48606_48668 (
    .I(net_48606),
    .O(net_48668)
  );
  InMux inmux_11_29_48616_48669 (
    .I(net_48616),
    .O(net_48669)
  );
  InMux inmux_11_30_48737_48766 (
    .I(net_48737),
    .O(net_48766)
  );
  InMux inmux_11_30_48737_48778 (
    .I(net_48737),
    .O(net_48778)
  );
  InMux inmux_11_30_48738_48767 (
    .I(net_48738),
    .O(net_48767)
  );
  InMux inmux_11_30_48738_48779 (
    .I(net_48738),
    .O(net_48779)
  );
  InMux inmux_11_30_48742_48768 (
    .I(net_48742),
    .O(net_48768)
  );
  InMux inmux_11_30_48742_48780 (
    .I(net_48742),
    .O(net_48780)
  );
  InMux inmux_11_30_48747_48765 (
    .I(net_48747),
    .O(net_48765)
  );
  InMux inmux_11_30_48747_48777 (
    .I(net_48747),
    .O(net_48777)
  );
  InMux inmux_11_7_45907_45933 (
    .I(net_45907),
    .O(net_45933)
  );
  CEMux inmux_11_7_45908_45976 (
    .I(net_45908),
    .O(net_45976)
  );
  InMux inmux_11_7_45911_45931 (
    .I(net_45911),
    .O(net_45931)
  );
  InMux inmux_11_7_45912_45932 (
    .I(net_45912),
    .O(net_45932)
  );
  InMux inmux_11_7_45921_45943 (
    .I(net_45921),
    .O(net_45943)
  );
  InMux inmux_11_7_45921_45974 (
    .I(net_45921),
    .O(net_45974)
  );
  InMux inmux_11_7_45923_45945 (
    .I(net_45923),
    .O(net_45945)
  );
  InMux inmux_11_7_45923_45972 (
    .I(net_45923),
    .O(net_45972)
  );
  InMux inmux_11_7_45924_45930 (
    .I(net_45924),
    .O(net_45930)
  );
  ClkMux inmux_11_7_5_45977 (
    .I(net_5),
    .O(net_45977)
  );
  InMux inmux_11_8_46020_46072 (
    .I(net_46020),
    .O(net_46072)
  );
  InMux inmux_11_8_46021_46078 (
    .I(net_46021),
    .O(net_46078)
  );
  InMux inmux_11_8_46022_46091 (
    .I(net_46022),
    .O(net_46091)
  );
  InMux inmux_11_8_46023_46066 (
    .I(net_46023),
    .O(net_46066)
  );
  InMux inmux_11_8_46024_46084 (
    .I(net_46024),
    .O(net_46084)
  );
  InMux inmux_11_8_46028_46054 (
    .I(net_46028),
    .O(net_46054)
  );
  InMux inmux_11_8_46030_46073 (
    .I(net_46030),
    .O(net_46073)
  );
  InMux inmux_11_8_46030_46085 (
    .I(net_46030),
    .O(net_46085)
  );
  InMux inmux_11_8_46030_46090 (
    .I(net_46030),
    .O(net_46090)
  );
  InMux inmux_11_8_46030_46097 (
    .I(net_46030),
    .O(net_46097)
  );
  InMux inmux_11_8_46034_46095 (
    .I(net_46034),
    .O(net_46095)
  );
  InMux inmux_11_8_46035_46060 (
    .I(net_46035),
    .O(net_46060)
  );
  InMux inmux_11_8_46035_46067 (
    .I(net_46035),
    .O(net_46067)
  );
  InMux inmux_11_8_46035_46079 (
    .I(net_46035),
    .O(net_46079)
  );
  InMux inmux_11_8_46037_46061 (
    .I(net_46037),
    .O(net_46061)
  );
  InMux inmux_11_8_46058_46068 (
    .I(net_46058),
    .O(net_46068)
  );
  InMux inmux_11_8_46064_46074 (
    .I(net_46064),
    .O(net_46074)
  );
  InMux inmux_11_8_46070_46080 (
    .I(net_46070),
    .O(net_46080)
  );
  InMux inmux_11_8_46076_46086 (
    .I(net_46076),
    .O(net_46086)
  );
  InMux inmux_11_8_46082_46092 (
    .I(net_46082),
    .O(net_46092)
  );
  InMux inmux_11_8_46088_46098 (
    .I(net_46088),
    .O(net_46098)
  );
  InMux inmux_11_9_46145_46212 (
    .I(net_46145),
    .O(net_46212)
  );
  InMux inmux_11_9_46146_46201 (
    .I(net_46146),
    .O(net_46201)
  );
  InMux inmux_11_9_46147_46207 (
    .I(net_46147),
    .O(net_46207)
  );
  InMux inmux_11_9_46148_46218 (
    .I(net_46148),
    .O(net_46218)
  );
  InMux inmux_11_9_46149_46200 (
    .I(net_46149),
    .O(net_46200)
  );
  InMux inmux_11_9_46149_46209 (
    .I(net_46149),
    .O(net_46209)
  );
  InMux inmux_11_9_46149_46214 (
    .I(net_46149),
    .O(net_46214)
  );
  InMux inmux_11_9_46150_46213 (
    .I(net_46150),
    .O(net_46213)
  );
  CEMux inmux_11_9_46154_46222 (
    .I(net_46154),
    .O(net_46222)
  );
  InMux inmux_11_9_46155_46179 (
    .I(net_46155),
    .O(net_46179)
  );
  InMux inmux_11_9_46155_46220 (
    .I(net_46155),
    .O(net_46220)
  );
  InMux inmux_11_9_46156_46183 (
    .I(net_46156),
    .O(net_46183)
  );
  InMux inmux_11_9_46156_46219 (
    .I(net_46156),
    .O(net_46219)
  );
  InMux inmux_11_9_46157_46203 (
    .I(net_46157),
    .O(net_46203)
  );
  InMux inmux_11_9_46157_46208 (
    .I(net_46157),
    .O(net_46208)
  );
  InMux inmux_11_9_46157_46215 (
    .I(net_46157),
    .O(net_46215)
  );
  InMux inmux_11_9_46158_46202 (
    .I(net_46158),
    .O(net_46202)
  );
  InMux inmux_11_9_46165_46197 (
    .I(net_46165),
    .O(net_46197)
  );
  InMux inmux_11_9_46165_46221 (
    .I(net_46165),
    .O(net_46221)
  );
  InMux inmux_11_9_46167_46206 (
    .I(net_46167),
    .O(net_46206)
  );
  ClkMux inmux_11_9_5_46223 (
    .I(net_5),
    .O(net_46223)
  );
  InMux inmux_12_11_50220_50260 (
    .I(net_50220),
    .O(net_50260)
  );
  InMux inmux_12_11_50220_50284 (
    .I(net_50220),
    .O(net_50284)
  );
  InMux inmux_12_11_50223_50261 (
    .I(net_50223),
    .O(net_50261)
  );
  InMux inmux_12_11_50226_50265 (
    .I(net_50226),
    .O(net_50265)
  );
  InMux inmux_12_11_50226_50272 (
    .I(net_50226),
    .O(net_50272)
  );
  InMux inmux_12_11_50227_50273 (
    .I(net_50227),
    .O(net_50273)
  );
  InMux inmux_12_11_50229_50253 (
    .I(net_50229),
    .O(net_50253)
  );
  InMux inmux_12_11_50230_50259 (
    .I(net_50230),
    .O(net_50259)
  );
  InMux inmux_12_11_50234_50292 (
    .I(net_50234),
    .O(net_50292)
  );
  InMux inmux_12_11_50239_50271 (
    .I(net_50239),
    .O(net_50271)
  );
  InMux inmux_12_11_50240_50262 (
    .I(net_50240),
    .O(net_50262)
  );
  InMux inmux_12_11_50240_50274 (
    .I(net_50240),
    .O(net_50274)
  );
  CEMux inmux_12_11_50247_50299 (
    .I(net_50247),
    .O(net_50299)
  );
  ClkMux inmux_12_11_5_50300 (
    .I(net_5),
    .O(net_50300)
  );
  InMux inmux_12_12_50343_50414 (
    .I(net_50343),
    .O(net_50414)
  );
  InMux inmux_12_12_50344_50384 (
    .I(net_50344),
    .O(net_50384)
  );
  InMux inmux_12_12_50345_50390 (
    .I(net_50345),
    .O(net_50390)
  );
  InMux inmux_12_12_50346_50389 (
    .I(net_50346),
    .O(net_50389)
  );
  InMux inmux_12_12_50347_50395 (
    .I(net_50347),
    .O(net_50395)
  );
  InMux inmux_12_12_50348_50413 (
    .I(net_50348),
    .O(net_50413)
  );
  InMux inmux_12_12_50349_50402 (
    .I(net_50349),
    .O(net_50402)
  );
  InMux inmux_12_12_50351_50420 (
    .I(net_50351),
    .O(net_50420)
  );
  InMux inmux_12_12_50353_50401 (
    .I(net_50353),
    .O(net_50401)
  );
  CEMux inmux_12_12_50354_50422 (
    .I(net_50354),
    .O(net_50422)
  );
  InMux inmux_12_12_50355_50408 (
    .I(net_50355),
    .O(net_50408)
  );
  InMux inmux_12_12_50356_50419 (
    .I(net_50356),
    .O(net_50419)
  );
  InMux inmux_12_12_50359_50378 (
    .I(net_50359),
    .O(net_50378)
  );
  InMux inmux_12_12_50360_50377 (
    .I(net_50360),
    .O(net_50377)
  );
  InMux inmux_12_12_50361_50383 (
    .I(net_50361),
    .O(net_50383)
  );
  InMux inmux_12_12_50370_50407 (
    .I(net_50370),
    .O(net_50407)
  );
  InMux inmux_12_12_50371_50396 (
    .I(net_50371),
    .O(net_50396)
  );
  InMux inmux_12_12_50375_50385 (
    .I(net_50375),
    .O(net_50385)
  );
  InMux inmux_12_12_50381_50391 (
    .I(net_50381),
    .O(net_50391)
  );
  InMux inmux_12_12_50387_50397 (
    .I(net_50387),
    .O(net_50397)
  );
  InMux inmux_12_12_50393_50403 (
    .I(net_50393),
    .O(net_50403)
  );
  InMux inmux_12_12_50399_50409 (
    .I(net_50399),
    .O(net_50409)
  );
  InMux inmux_12_12_50405_50415 (
    .I(net_50405),
    .O(net_50415)
  );
  InMux inmux_12_12_50411_50421 (
    .I(net_50411),
    .O(net_50421)
  );
  ClkMux inmux_12_12_5_50423 (
    .I(net_5),
    .O(net_50423)
  );
  InMux inmux_12_13_50461_50502 (
    .I(net_50461),
    .O(net_50502)
  );
  InMux inmux_12_13_50466_50518 (
    .I(net_50466),
    .O(net_50518)
  );
  InMux inmux_12_13_50467_50536 (
    .I(net_50467),
    .O(net_50536)
  );
  InMux inmux_12_13_50468_50525 (
    .I(net_50468),
    .O(net_50525)
  );
  InMux inmux_12_13_50469_50524 (
    .I(net_50469),
    .O(net_50524)
  );
  InMux inmux_12_13_50471_50543 (
    .I(net_50471),
    .O(net_50543)
  );
  InMux inmux_12_13_50474_50507 (
    .I(net_50474),
    .O(net_50507)
  );
  InMux inmux_12_13_50475_50537 (
    .I(net_50475),
    .O(net_50537)
  );
  InMux inmux_12_13_50477_50513 (
    .I(net_50477),
    .O(net_50513)
  );
  InMux inmux_12_13_50478_50512 (
    .I(net_50478),
    .O(net_50512)
  );
  InMux inmux_12_13_50479_50542 (
    .I(net_50479),
    .O(net_50542)
  );
  InMux inmux_12_13_50481_50530 (
    .I(net_50481),
    .O(net_50530)
  );
  InMux inmux_12_13_50483_50500 (
    .I(net_50483),
    .O(net_50500)
  );
  InMux inmux_12_13_50484_50501 (
    .I(net_50484),
    .O(net_50501)
  );
  InMux inmux_12_13_50485_50519 (
    .I(net_50485),
    .O(net_50519)
  );
  InMux inmux_12_13_50492_50531 (
    .I(net_50492),
    .O(net_50531)
  );
  CEMux inmux_12_13_50493_50545 (
    .I(net_50493),
    .O(net_50545)
  );
  InMux inmux_12_13_50495_50506 (
    .I(net_50495),
    .O(net_50506)
  );
  InMux inmux_12_13_50498_50508 (
    .I(net_50498),
    .O(net_50508)
  );
  InMux inmux_12_13_50504_50514 (
    .I(net_50504),
    .O(net_50514)
  );
  InMux inmux_12_13_50510_50520 (
    .I(net_50510),
    .O(net_50520)
  );
  InMux inmux_12_13_50516_50526 (
    .I(net_50516),
    .O(net_50526)
  );
  InMux inmux_12_13_50522_50532 (
    .I(net_50522),
    .O(net_50532)
  );
  InMux inmux_12_13_50528_50538 (
    .I(net_50528),
    .O(net_50538)
  );
  InMux inmux_12_13_50534_50544 (
    .I(net_50534),
    .O(net_50544)
  );
  ClkMux inmux_12_13_5_50546 (
    .I(net_5),
    .O(net_50546)
  );
  InMux inmux_12_14_50593_50622 (
    .I(net_50593),
    .O(net_50622)
  );
  InMux inmux_12_14_50597_50666 (
    .I(net_50597),
    .O(net_50666)
  );
  InMux inmux_12_14_50598_50634 (
    .I(net_50598),
    .O(net_50634)
  );
  InMux inmux_12_14_50598_50667 (
    .I(net_50598),
    .O(net_50667)
  );
  InMux inmux_12_14_50599_50623 (
    .I(net_50599),
    .O(net_50623)
  );
  InMux inmux_12_14_50600_50665 (
    .I(net_50600),
    .O(net_50665)
  );
  InMux inmux_12_14_50601_50635 (
    .I(net_50601),
    .O(net_50635)
  );
  InMux inmux_12_14_50601_50640 (
    .I(net_50601),
    .O(net_50640)
  );
  InMux inmux_12_14_50602_50624 (
    .I(net_50602),
    .O(net_50624)
  );
  InMux inmux_12_14_50603_50649 (
    .I(net_50603),
    .O(net_50649)
  );
  InMux inmux_12_14_50609_50636 (
    .I(net_50609),
    .O(net_50636)
  );
  InMux inmux_12_14_50613_50664 (
    .I(net_50613),
    .O(net_50664)
  );
  InMux inmux_12_14_50615_50637 (
    .I(net_50615),
    .O(net_50637)
  );
  CEMux inmux_12_14_50616_50668 (
    .I(net_50616),
    .O(net_50668)
  );
  InMux inmux_12_14_50617_50654 (
    .I(net_50617),
    .O(net_50654)
  );
  InMux inmux_12_14_50620_50631 (
    .I(net_50620),
    .O(net_50631)
  );
  ClkMux inmux_12_14_5_50669 (
    .I(net_5),
    .O(net_50669)
  );
  InMux inmux_12_15_50712_50745 (
    .I(net_50712),
    .O(net_50745)
  );
  InMux inmux_12_15_50713_50770 (
    .I(net_50713),
    .O(net_50770)
  );
  InMux inmux_12_15_50713_50777 (
    .I(net_50713),
    .O(net_50777)
  );
  InMux inmux_12_15_50716_50757 (
    .I(net_50716),
    .O(net_50757)
  );
  InMux inmux_12_15_50718_50752 (
    .I(net_50718),
    .O(net_50752)
  );
  InMux inmux_12_15_50718_50769 (
    .I(net_50718),
    .O(net_50769)
  );
  InMux inmux_12_15_50722_50760 (
    .I(net_50722),
    .O(net_50760)
  );
  InMux inmux_12_15_50722_50763 (
    .I(net_50722),
    .O(net_50763)
  );
  InMux inmux_12_15_50724_50775 (
    .I(net_50724),
    .O(net_50775)
  );
  InMux inmux_12_15_50726_50789 (
    .I(net_50726),
    .O(net_50789)
  );
  InMux inmux_12_15_50728_50778 (
    .I(net_50728),
    .O(net_50778)
  );
  InMux inmux_12_15_50735_50772 (
    .I(net_50735),
    .O(net_50772)
  );
  InMux inmux_12_15_50740_50758 (
    .I(net_50740),
    .O(net_50758)
  );
  InMux inmux_12_15_50743_50759 (
    .I(net_50743),
    .O(net_50759)
  );
  InMux inmux_12_15_50743_50771 (
    .I(net_50743),
    .O(net_50771)
  );
  InMux inmux_12_15_50743_50776 (
    .I(net_50743),
    .O(net_50776)
  );
  ClkMux inmux_12_15_5_50792 (
    .I(net_5),
    .O(net_50792)
  );
  CEMux inmux_12_15_6_50791 (
    .I(net_6),
    .O(net_50791)
  );
  InMux inmux_12_16_50835_50899 (
    .I(net_50835),
    .O(net_50899)
  );
  InMux inmux_12_16_50835_50906 (
    .I(net_50835),
    .O(net_50906)
  );
  InMux inmux_12_16_50836_50898 (
    .I(net_50836),
    .O(net_50898)
  );
  InMux inmux_12_16_50854_50883 (
    .I(net_50854),
    .O(net_50883)
  );
  InMux inmux_12_16_50861_50876 (
    .I(net_50861),
    .O(net_50876)
  );
  InMux inmux_12_16_50861_50905 (
    .I(net_50861),
    .O(net_50905)
  );
  CEMux inmux_12_16_50862_50914 (
    .I(net_50862),
    .O(net_50914)
  );
  InMux inmux_12_16_50865_50893 (
    .I(net_50865),
    .O(net_50893)
  );
  ClkMux inmux_12_16_5_50915 (
    .I(net_5),
    .O(net_50915)
  );
  CEMux inmux_12_17_50960_51037 (
    .I(net_50960),
    .O(net_51037)
  );
  InMux inmux_12_17_50962_51012 (
    .I(net_50962),
    .O(net_51012)
  );
  InMux inmux_12_17_50963_50999 (
    .I(net_50963),
    .O(net_50999)
  );
  InMux inmux_12_17_50967_50993 (
    .I(net_50967),
    .O(net_50993)
  );
  InMux inmux_12_17_50971_51027 (
    .I(net_50971),
    .O(net_51027)
  );
  InMux inmux_12_17_50980_51022 (
    .I(net_50980),
    .O(net_51022)
  );
  ClkMux inmux_12_17_5_51038 (
    .I(net_5),
    .O(net_51038)
  );
  InMux inmux_12_18_51082_51127 (
    .I(net_51082),
    .O(net_51127)
  );
  InMux inmux_12_18_51085_51128 (
    .I(net_51085),
    .O(net_51128)
  );
  InMux inmux_12_18_51086_51129 (
    .I(net_51086),
    .O(net_51129)
  );
  InMux inmux_12_18_51088_51117 (
    .I(net_51088),
    .O(net_51117)
  );
  InMux inmux_12_18_51095_51115 (
    .I(net_51095),
    .O(net_51115)
  );
  InMux inmux_12_18_51099_51116 (
    .I(net_51099),
    .O(net_51116)
  );
  InMux inmux_12_18_51101_51114 (
    .I(net_51101),
    .O(net_51114)
  );
  InMux inmux_12_18_51103_51157 (
    .I(net_51103),
    .O(net_51157)
  );
  InMux inmux_12_18_51105_51144 (
    .I(net_51105),
    .O(net_51144)
  );
  InMux inmux_12_18_51106_51126 (
    .I(net_51106),
    .O(net_51126)
  );
  ClkMux inmux_12_18_5_51161 (
    .I(net_5),
    .O(net_51161)
  );
  CEMux inmux_12_18_6_51160 (
    .I(net_6),
    .O(net_51160)
  );
  InMux inmux_12_19_51210_51261 (
    .I(net_51210),
    .O(net_51261)
  );
  InMux inmux_12_19_51213_51251 (
    .I(net_51213),
    .O(net_51251)
  );
  InMux inmux_12_19_51214_51250 (
    .I(net_51214),
    .O(net_51250)
  );
  InMux inmux_12_19_51215_51263 (
    .I(net_51215),
    .O(net_51263)
  );
  InMux inmux_12_19_51215_51282 (
    .I(net_51215),
    .O(net_51282)
  );
  InMux inmux_12_19_51216_51252 (
    .I(net_51216),
    .O(net_51252)
  );
  InMux inmux_12_19_51220_51256 (
    .I(net_51220),
    .O(net_51256)
  );
  CEMux inmux_12_19_51222_51283 (
    .I(net_51222),
    .O(net_51283)
  );
  InMux inmux_12_19_51228_51276 (
    .I(net_51228),
    .O(net_51276)
  );
  InMux inmux_12_19_51231_51280 (
    .I(net_51231),
    .O(net_51280)
  );
  InMux inmux_12_19_51235_51249 (
    .I(net_51235),
    .O(net_51249)
  );
  ClkMux inmux_12_19_5_51284 (
    .I(net_5),
    .O(net_51284)
  );
  InMux inmux_12_20_51343_51367 (
    .I(net_51343),
    .O(net_51367)
  );
  ClkMux inmux_12_20_5_51407 (
    .I(net_5),
    .O(net_51407)
  );
  CEMux inmux_12_20_8_51406 (
    .I(net_8),
    .O(net_51406)
  );
  InMux inmux_12_21_51452_51528 (
    .I(net_51452),
    .O(net_51528)
  );
  InMux inmux_12_21_51456_51526 (
    .I(net_51456),
    .O(net_51526)
  );
  InMux inmux_12_21_51460_51527 (
    .I(net_51460),
    .O(net_51527)
  );
  CEMux inmux_12_21_51461_51529 (
    .I(net_51461),
    .O(net_51529)
  );
  SRMux inmux_12_21_51470_51531 (
    .I(net_51470),
    .O(net_51531)
  );
  InMux inmux_12_21_51471_51484 (
    .I(net_51471),
    .O(net_51484)
  );
  InMux inmux_12_21_51471_51510 (
    .I(net_51471),
    .O(net_51510)
  );
  InMux inmux_12_21_51471_51525 (
    .I(net_51471),
    .O(net_51525)
  );
  InMux inmux_12_21_51473_51498 (
    .I(net_51473),
    .O(net_51498)
  );
  InMux inmux_12_21_51473_51508 (
    .I(net_51473),
    .O(net_51508)
  );
  InMux inmux_12_21_51473_51522 (
    .I(net_51473),
    .O(net_51522)
  );
  InMux inmux_12_21_51477_51485 (
    .I(net_51477),
    .O(net_51485)
  );
  InMux inmux_12_21_51477_51521 (
    .I(net_51477),
    .O(net_51521)
  );
  ClkMux inmux_12_21_5_51530 (
    .I(net_5),
    .O(net_51530)
  );
  InMux inmux_12_23_51719_51730 (
    .I(net_51719),
    .O(net_51730)
  );
  ClkMux inmux_12_23_5_51776 (
    .I(net_5),
    .O(net_51776)
  );
  InMux inmux_12_27_52195_52234 (
    .I(net_52195),
    .O(net_52234)
  );
  InMux inmux_12_27_52197_52223 (
    .I(net_52197),
    .O(net_52223)
  );
  CEMux inmux_12_27_52199_52267 (
    .I(net_52199),
    .O(net_52267)
  );
  InMux inmux_12_27_52206_52266 (
    .I(net_52206),
    .O(net_52266)
  );
  InMux inmux_12_27_52207_52258 (
    .I(net_52207),
    .O(net_52258)
  );
  InMux inmux_12_27_52208_52252 (
    .I(net_52208),
    .O(net_52252)
  );
  InMux inmux_12_27_52209_52229 (
    .I(net_52209),
    .O(net_52229)
  );
  InMux inmux_12_27_52211_52246 (
    .I(net_52211),
    .O(net_52246)
  );
  InMux inmux_12_27_52215_52257 (
    .I(net_52215),
    .O(net_52257)
  );
  InMux inmux_12_27_52215_52264 (
    .I(net_52215),
    .O(net_52264)
  );
  InMux inmux_12_27_52218_52241 (
    .I(net_52218),
    .O(net_52241)
  );
  InMux inmux_12_27_52226_52236 (
    .I(net_52226),
    .O(net_52236)
  );
  InMux inmux_12_27_52232_52242 (
    .I(net_52232),
    .O(net_52242)
  );
  InMux inmux_12_27_52238_52248 (
    .I(net_52238),
    .O(net_52248)
  );
  InMux inmux_12_27_52244_52254 (
    .I(net_52244),
    .O(net_52254)
  );
  ClkMux inmux_12_27_5_52268 (
    .I(net_5),
    .O(net_52268)
  );
  CEMux inmux_12_28_52313_52390 (
    .I(net_52313),
    .O(net_52390)
  );
  InMux inmux_12_28_52320_52356 (
    .I(net_52320),
    .O(net_52356)
  );
  InMux inmux_12_28_52321_52352 (
    .I(net_52321),
    .O(net_52352)
  );
  InMux inmux_12_28_52322_52353 (
    .I(net_52322),
    .O(net_52353)
  );
  InMux inmux_12_28_52336_52358 (
    .I(net_52336),
    .O(net_52358)
  );
  ClkMux inmux_12_28_5_52391 (
    .I(net_5),
    .O(net_52391)
  );
  CEMux inmux_12_8_49862_49930 (
    .I(net_49862),
    .O(net_49930)
  );
  InMux inmux_12_8_49866_49922 (
    .I(net_49866),
    .O(net_49922)
  );
  InMux inmux_12_8_49872_49892 (
    .I(net_49872),
    .O(net_49892)
  );
  InMux inmux_12_8_49875_49923 (
    .I(net_49875),
    .O(net_49923)
  );
  InMux inmux_12_8_49876_49915 (
    .I(net_49876),
    .O(net_49915)
  );
  InMux inmux_12_8_49880_49920 (
    .I(net_49880),
    .O(net_49920)
  );
  ClkMux inmux_12_8_5_49931 (
    .I(net_5),
    .O(net_49931)
  );
  InMux inmux_13_11_54064_54120 (
    .I(net_54064),
    .O(net_54120)
  );
  CEMux inmux_13_11_54069_54130 (
    .I(net_54069),
    .O(net_54130)
  );
  InMux inmux_13_11_54081_54090 (
    .I(net_54081),
    .O(net_54090)
  );
  ClkMux inmux_13_11_5_54131 (
    .I(net_5),
    .O(net_54131)
  );
  InMux inmux_13_12_54175_54227 (
    .I(net_54175),
    .O(net_54227)
  );
  CEMux inmux_13_12_54176_54253 (
    .I(net_54176),
    .O(net_54253)
  );
  InMux inmux_13_12_54177_54222 (
    .I(net_54177),
    .O(net_54222)
  );
  InMux inmux_13_12_54178_54252 (
    .I(net_54178),
    .O(net_54252)
  );
  InMux inmux_13_12_54179_54210 (
    .I(net_54179),
    .O(net_54210)
  );
  InMux inmux_13_12_54179_54234 (
    .I(net_54179),
    .O(net_54234)
  );
  InMux inmux_13_12_54186_54246 (
    .I(net_54186),
    .O(net_54246)
  );
  InMux inmux_13_12_54187_54209 (
    .I(net_54187),
    .O(net_54209)
  );
  InMux inmux_13_12_54187_54219 (
    .I(net_54187),
    .O(net_54219)
  );
  InMux inmux_13_12_54187_54228 (
    .I(net_54187),
    .O(net_54228)
  );
  InMux inmux_13_12_54187_54245 (
    .I(net_54187),
    .O(net_54245)
  );
  InMux inmux_13_12_54188_54225 (
    .I(net_54188),
    .O(net_54225)
  );
  InMux inmux_13_12_54189_54214 (
    .I(net_54189),
    .O(net_54214)
  );
  InMux inmux_13_12_54190_54207 (
    .I(net_54190),
    .O(net_54207)
  );
  InMux inmux_13_12_54190_54221 (
    .I(net_54190),
    .O(net_54221)
  );
  InMux inmux_13_12_54190_54226 (
    .I(net_54190),
    .O(net_54226)
  );
  InMux inmux_13_12_54190_54243 (
    .I(net_54190),
    .O(net_54243)
  );
  InMux inmux_13_12_54191_54215 (
    .I(net_54191),
    .O(net_54215)
  );
  InMux inmux_13_12_54193_54220 (
    .I(net_54193),
    .O(net_54220)
  );
  InMux inmux_13_12_54195_54244 (
    .I(net_54195),
    .O(net_54244)
  );
  InMux inmux_13_12_54202_54208 (
    .I(net_54202),
    .O(net_54208)
  );
  InMux inmux_13_12_54205_54238 (
    .I(net_54205),
    .O(net_54238)
  );
  ClkMux inmux_13_12_5_54254 (
    .I(net_5),
    .O(net_54254)
  );
  InMux inmux_13_13_54297_54349 (
    .I(net_54297),
    .O(net_54349)
  );
  InMux inmux_13_13_54299_54332 (
    .I(net_54299),
    .O(net_54332)
  );
  InMux inmux_13_13_54300_54333 (
    .I(net_54300),
    .O(net_54333)
  );
  InMux inmux_13_13_54302_54343 (
    .I(net_54302),
    .O(net_54343)
  );
  InMux inmux_13_13_54302_54374 (
    .I(net_54302),
    .O(net_54374)
  );
  InMux inmux_13_13_54305_54345 (
    .I(net_54305),
    .O(net_54345)
  );
  InMux inmux_13_13_54308_54373 (
    .I(net_54308),
    .O(net_54373)
  );
  InMux inmux_13_13_54309_54331 (
    .I(net_54309),
    .O(net_54331)
  );
  InMux inmux_13_13_54310_54330 (
    .I(net_54310),
    .O(net_54330)
  );
  InMux inmux_13_13_54312_54344 (
    .I(net_54312),
    .O(net_54344)
  );
  InMux inmux_13_13_54312_54375 (
    .I(net_54312),
    .O(net_54375)
  );
  InMux inmux_13_13_54316_54372 (
    .I(net_54316),
    .O(net_54372)
  );
  InMux inmux_13_13_54318_54338 (
    .I(net_54318),
    .O(net_54338)
  );
  InMux inmux_13_13_54319_54356 (
    .I(net_54319),
    .O(net_54356)
  );
  InMux inmux_13_13_54323_54369 (
    .I(net_54323),
    .O(net_54369)
  );
  InMux inmux_13_13_54325_54348 (
    .I(net_54325),
    .O(net_54348)
  );
  InMux inmux_13_13_54326_54342 (
    .I(net_54326),
    .O(net_54342)
  );
  InMux inmux_13_13_54328_54363 (
    .I(net_54328),
    .O(net_54363)
  );
  ClkMux inmux_13_13_5_54377 (
    .I(net_5),
    .O(net_54377)
  );
  CEMux inmux_13_13_6_54376 (
    .I(net_6),
    .O(net_54376)
  );
  InMux inmux_13_14_54426_54472 (
    .I(net_54426),
    .O(net_54472)
  );
  InMux inmux_13_14_54427_54480 (
    .I(net_54427),
    .O(net_54480)
  );
  InMux inmux_13_14_54428_54473 (
    .I(net_54428),
    .O(net_54473)
  );
  InMux inmux_13_14_54428_54490 (
    .I(net_54428),
    .O(net_54490)
  );
  CEMux inmux_13_14_54431_54499 (
    .I(net_54431),
    .O(net_54499)
  );
  InMux inmux_13_14_54433_54491 (
    .I(net_54433),
    .O(net_54491)
  );
  InMux inmux_13_14_54434_54456 (
    .I(net_54434),
    .O(net_54456)
  );
  InMux inmux_13_14_54435_54453 (
    .I(net_54435),
    .O(net_54453)
  );
  InMux inmux_13_14_54437_54483 (
    .I(net_54437),
    .O(net_54483)
  );
  InMux inmux_13_14_54442_54455 (
    .I(net_54442),
    .O(net_54455)
  );
  InMux inmux_13_14_54444_54454 (
    .I(net_54444),
    .O(net_54454)
  );
  InMux inmux_13_14_54444_54471 (
    .I(net_54444),
    .O(net_54471)
  );
  InMux inmux_13_14_54444_54492 (
    .I(net_54444),
    .O(net_54492)
  );
  InMux inmux_13_14_54446_54459 (
    .I(net_54446),
    .O(net_54459)
  );
  InMux inmux_13_14_54446_54478 (
    .I(net_54446),
    .O(net_54478)
  );
  InMux inmux_13_14_54447_54496 (
    .I(net_54447),
    .O(net_54496)
  );
  InMux inmux_13_14_54449_54467 (
    .I(net_54449),
    .O(net_54467)
  );
  InMux inmux_13_14_54449_54474 (
    .I(net_54449),
    .O(net_54474)
  );
  InMux inmux_13_14_54450_54461 (
    .I(net_54450),
    .O(net_54461)
  );
  InMux inmux_13_14_54451_54489 (
    .I(net_54451),
    .O(net_54489)
  );
  ClkMux inmux_13_14_5_54500 (
    .I(net_5),
    .O(net_54500)
  );
  InMux inmux_13_15_54545_54609 (
    .I(net_54545),
    .O(net_54609)
  );
  InMux inmux_13_15_54548_54618 (
    .I(net_54548),
    .O(net_54618)
  );
  InMux inmux_13_15_54553_54620 (
    .I(net_54553),
    .O(net_54620)
  );
  InMux inmux_13_15_54555_54579 (
    .I(net_54555),
    .O(net_54579)
  );
  InMux inmux_13_15_54559_54595 (
    .I(net_54559),
    .O(net_54595)
  );
  InMux inmux_13_15_54560_54577 (
    .I(net_54560),
    .O(net_54577)
  );
  InMux inmux_13_15_54561_54614 (
    .I(net_54561),
    .O(net_54614)
  );
  InMux inmux_13_15_54562_54582 (
    .I(net_54562),
    .O(net_54582)
  );
  InMux inmux_13_15_54564_54589 (
    .I(net_54564),
    .O(net_54589)
  );
  InMux inmux_13_15_54565_54576 (
    .I(net_54565),
    .O(net_54576)
  );
  InMux inmux_13_15_54569_54596 (
    .I(net_54569),
    .O(net_54596)
  );
  InMux inmux_13_15_54570_54578 (
    .I(net_54570),
    .O(net_54578)
  );
  InMux inmux_13_15_54570_54621 (
    .I(net_54570),
    .O(net_54621)
  );
  InMux inmux_13_15_54572_54619 (
    .I(net_54572),
    .O(net_54619)
  );
  InMux inmux_13_15_54573_54603 (
    .I(net_54573),
    .O(net_54603)
  );
  ClkMux inmux_13_15_5_54623 (
    .I(net_5),
    .O(net_54623)
  );
  CEMux inmux_13_15_8_54622 (
    .I(net_8),
    .O(net_54622)
  );
  InMux inmux_13_16_54668_54718 (
    .I(net_54668),
    .O(net_54718)
  );
  InMux inmux_13_16_54670_54713 (
    .I(net_54670),
    .O(net_54713)
  );
  InMux inmux_13_16_54672_54701 (
    .I(net_54672),
    .O(net_54701)
  );
  CEMux inmux_13_16_54677_54745 (
    .I(net_54677),
    .O(net_54745)
  );
  InMux inmux_13_16_54680_54724 (
    .I(net_54680),
    .O(net_54724)
  );
  InMux inmux_13_16_54682_54742 (
    .I(net_54682),
    .O(net_54742)
  );
  InMux inmux_13_16_54685_54700 (
    .I(net_54685),
    .O(net_54700)
  );
  InMux inmux_13_16_54686_54706 (
    .I(net_54686),
    .O(net_54706)
  );
  InMux inmux_13_16_54687_54736 (
    .I(net_54687),
    .O(net_54736)
  );
  InMux inmux_13_16_54689_54707 (
    .I(net_54689),
    .O(net_54707)
  );
  InMux inmux_13_16_54690_54719 (
    .I(net_54690),
    .O(net_54719)
  );
  InMux inmux_13_16_54692_54712 (
    .I(net_54692),
    .O(net_54712)
  );
  InMux inmux_13_16_54693_54737 (
    .I(net_54693),
    .O(net_54737)
  );
  InMux inmux_13_16_54694_54743 (
    .I(net_54694),
    .O(net_54743)
  );
  InMux inmux_13_16_54695_54730 (
    .I(net_54695),
    .O(net_54730)
  );
  InMux inmux_13_16_54696_54731 (
    .I(net_54696),
    .O(net_54731)
  );
  InMux inmux_13_16_54697_54725 (
    .I(net_54697),
    .O(net_54725)
  );
  InMux inmux_13_16_54698_54708 (
    .I(net_54698),
    .O(net_54708)
  );
  InMux inmux_13_16_54704_54714 (
    .I(net_54704),
    .O(net_54714)
  );
  InMux inmux_13_16_54710_54720 (
    .I(net_54710),
    .O(net_54720)
  );
  InMux inmux_13_16_54716_54726 (
    .I(net_54716),
    .O(net_54726)
  );
  InMux inmux_13_16_54722_54732 (
    .I(net_54722),
    .O(net_54732)
  );
  InMux inmux_13_16_54728_54738 (
    .I(net_54728),
    .O(net_54738)
  );
  InMux inmux_13_16_54734_54744 (
    .I(net_54734),
    .O(net_54744)
  );
  ClkMux inmux_13_16_5_54746 (
    .I(net_5),
    .O(net_54746)
  );
  InMux inmux_13_17_54784_54825 (
    .I(net_54784),
    .O(net_54825)
  );
  InMux inmux_13_17_54789_54829 (
    .I(net_54789),
    .O(net_54829)
  );
  InMux inmux_13_17_54792_54854 (
    .I(net_54792),
    .O(net_54854)
  );
  InMux inmux_13_17_54793_54836 (
    .I(net_54793),
    .O(net_54836)
  );
  InMux inmux_13_17_54795_54824 (
    .I(net_54795),
    .O(net_54824)
  );
  InMux inmux_13_17_54797_54866 (
    .I(net_54797),
    .O(net_54866)
  );
  InMux inmux_13_17_54801_54835 (
    .I(net_54801),
    .O(net_54835)
  );
  InMux inmux_13_17_54803_54823 (
    .I(net_54803),
    .O(net_54823)
  );
  InMux inmux_13_17_54805_54865 (
    .I(net_54805),
    .O(net_54865)
  );
  InMux inmux_13_17_54806_54847 (
    .I(net_54806),
    .O(net_54847)
  );
  InMux inmux_13_17_54808_54842 (
    .I(net_54808),
    .O(net_54842)
  );
  InMux inmux_13_17_54811_54860 (
    .I(net_54811),
    .O(net_54860)
  );
  InMux inmux_13_17_54812_54859 (
    .I(net_54812),
    .O(net_54859)
  );
  InMux inmux_13_17_54814_54841 (
    .I(net_54814),
    .O(net_54841)
  );
  InMux inmux_13_17_54815_54830 (
    .I(net_54815),
    .O(net_54830)
  );
  CEMux inmux_13_17_54816_54868 (
    .I(net_54816),
    .O(net_54868)
  );
  InMux inmux_13_17_54818_54853 (
    .I(net_54818),
    .O(net_54853)
  );
  InMux inmux_13_17_54820_54848 (
    .I(net_54820),
    .O(net_54848)
  );
  InMux inmux_13_17_54821_54831 (
    .I(net_54821),
    .O(net_54831)
  );
  InMux inmux_13_17_54827_54837 (
    .I(net_54827),
    .O(net_54837)
  );
  InMux inmux_13_17_54833_54843 (
    .I(net_54833),
    .O(net_54843)
  );
  InMux inmux_13_17_54839_54849 (
    .I(net_54839),
    .O(net_54849)
  );
  InMux inmux_13_17_54845_54855 (
    .I(net_54845),
    .O(net_54855)
  );
  InMux inmux_13_17_54851_54861 (
    .I(net_54851),
    .O(net_54861)
  );
  InMux inmux_13_17_54857_54867 (
    .I(net_54857),
    .O(net_54867)
  );
  ClkMux inmux_13_17_5_54869 (
    .I(net_5),
    .O(net_54869)
  );
  InMux inmux_13_18_54912_54976 (
    .I(net_54912),
    .O(net_54976)
  );
  InMux inmux_13_18_54933_54970 (
    .I(net_54933),
    .O(net_54970)
  );
  InMux inmux_13_18_54943_54964 (
    .I(net_54943),
    .O(net_54964)
  );
  ClkMux inmux_13_18_5_54992 (
    .I(net_5),
    .O(net_54992)
  );
  CEMux inmux_13_18_8_54991 (
    .I(net_8),
    .O(net_54991)
  );
  InMux inmux_13_19_55042_55095 (
    .I(net_55042),
    .O(net_55095)
  );
  InMux inmux_13_19_55043_55107 (
    .I(net_55043),
    .O(net_55107)
  );
  InMux inmux_13_19_55049_55074 (
    .I(net_55049),
    .O(net_55074)
  );
  InMux inmux_13_19_55050_55075 (
    .I(net_55050),
    .O(net_55075)
  );
  InMux inmux_13_19_55052_55112 (
    .I(net_55052),
    .O(net_55112)
  );
  InMux inmux_13_19_55053_55092 (
    .I(net_55053),
    .O(net_55092)
  );
  InMux inmux_13_19_55055_55077 (
    .I(net_55055),
    .O(net_55077)
  );
  InMux inmux_13_19_55056_55105 (
    .I(net_55056),
    .O(net_55105)
  );
  InMux inmux_13_19_55057_55094 (
    .I(net_55057),
    .O(net_55094)
  );
  InMux inmux_13_19_55058_55076 (
    .I(net_55058),
    .O(net_55076)
  );
  InMux inmux_13_19_55062_55106 (
    .I(net_55062),
    .O(net_55106)
  );
  InMux inmux_13_19_55063_55093 (
    .I(net_55063),
    .O(net_55093)
  );
  InMux inmux_13_19_55064_55082 (
    .I(net_55064),
    .O(net_55082)
  );
  InMux inmux_13_19_55066_55104 (
    .I(net_55066),
    .O(net_55104)
  );
  ClkMux inmux_13_19_5_55115 (
    .I(net_5),
    .O(net_55115)
  );
  CEMux inmux_13_19_8_55114 (
    .I(net_8),
    .O(net_55114)
  );
  CEMux inmux_13_20_55169_55237 (
    .I(net_55169),
    .O(net_55237)
  );
  InMux inmux_13_20_55171_55234 (
    .I(net_55171),
    .O(net_55234)
  );
  InMux inmux_13_20_55172_55228 (
    .I(net_55172),
    .O(net_55228)
  );
  InMux inmux_13_20_55172_55235 (
    .I(net_55172),
    .O(net_55235)
  );
  InMux inmux_13_20_55175_55230 (
    .I(net_55175),
    .O(net_55230)
  );
  InMux inmux_13_20_55176_55227 (
    .I(net_55176),
    .O(net_55227)
  );
  InMux inmux_13_20_55176_55236 (
    .I(net_55176),
    .O(net_55236)
  );
  InMux inmux_13_20_55178_55229 (
    .I(net_55178),
    .O(net_55229)
  );
  InMux inmux_13_20_55181_55223 (
    .I(net_55181),
    .O(net_55223)
  );
  InMux inmux_13_20_55182_55194 (
    .I(net_55182),
    .O(net_55194)
  );
  InMux inmux_13_20_55183_55200 (
    .I(net_55183),
    .O(net_55200)
  );
  InMux inmux_13_20_55186_55233 (
    .I(net_55186),
    .O(net_55233)
  );
  InMux inmux_13_20_55187_55217 (
    .I(net_55187),
    .O(net_55217)
  );
  InMux inmux_13_20_55189_55212 (
    .I(net_55189),
    .O(net_55212)
  );
  ClkMux inmux_13_20_5_55238 (
    .I(net_5),
    .O(net_55238)
  );
  InMux inmux_13_21_55309_55351 (
    .I(net_55309),
    .O(net_55351)
  );
  InMux inmux_13_22_55405_55457 (
    .I(net_55405),
    .O(net_55457)
  );
  InMux inmux_13_22_55405_55481 (
    .I(net_55405),
    .O(net_55481)
  );
  InMux inmux_13_22_55417_55456 (
    .I(net_55417),
    .O(net_55456)
  );
  InMux inmux_13_22_55417_55480 (
    .I(net_55417),
    .O(net_55480)
  );
  InMux inmux_13_22_55418_55443 (
    .I(net_55418),
    .O(net_55443)
  );
  CEMux inmux_13_22_55422_55483 (
    .I(net_55422),
    .O(net_55483)
  );
  InMux inmux_13_22_55423_55455 (
    .I(net_55423),
    .O(net_55455)
  );
  InMux inmux_13_22_55423_55479 (
    .I(net_55423),
    .O(net_55479)
  );
  InMux inmux_13_22_55433_55458 (
    .I(net_55433),
    .O(net_55458)
  );
  InMux inmux_13_22_55433_55470 (
    .I(net_55433),
    .O(net_55470)
  );
  InMux inmux_13_22_55433_55482 (
    .I(net_55433),
    .O(net_55482)
  );
  ClkMux inmux_13_22_5_55484 (
    .I(net_5),
    .O(net_55484)
  );
  CEMux inmux_13_27_56021_56098 (
    .I(net_56021),
    .O(net_56098)
  );
  InMux inmux_13_27_56024_56079 (
    .I(net_56024),
    .O(net_56079)
  );
  InMux inmux_13_27_56025_56064 (
    .I(net_56025),
    .O(net_56064)
  );
  InMux inmux_13_27_56026_56067 (
    .I(net_56026),
    .O(net_56067)
  );
  InMux inmux_13_27_56030_56076 (
    .I(net_56030),
    .O(net_56076)
  );
  InMux inmux_13_27_56030_56085 (
    .I(net_56030),
    .O(net_56085)
  );
  InMux inmux_13_27_56030_56088 (
    .I(net_56030),
    .O(net_56088)
  );
  InMux inmux_13_27_56030_56095 (
    .I(net_56030),
    .O(net_56095)
  );
  InMux inmux_13_27_56031_56094 (
    .I(net_56031),
    .O(net_56094)
  );
  InMux inmux_13_27_56034_56066 (
    .I(net_56034),
    .O(net_56066)
  );
  InMux inmux_13_27_56036_56082 (
    .I(net_56036),
    .O(net_56082)
  );
  InMux inmux_13_27_56036_56091 (
    .I(net_56036),
    .O(net_56091)
  );
  InMux inmux_13_27_56037_56090 (
    .I(net_56037),
    .O(net_56090)
  );
  InMux inmux_13_27_56040_56084 (
    .I(net_56040),
    .O(net_56084)
  );
  InMux inmux_13_27_56040_56089 (
    .I(net_56040),
    .O(net_56089)
  );
  InMux inmux_13_27_56047_56065 (
    .I(net_56047),
    .O(net_56065)
  );
  ClkMux inmux_13_27_5_56099 (
    .I(net_5),
    .O(net_56099)
  );
  CEMux inmux_13_31_56534_56521 (
    .I(net_56534),
    .O(net_56521)
  );
  IoInMux inmux_13_31_56535_56515 (
    .I(net_56535),
    .O(net_56515)
  );
  ClkMux inmux_13_31_5_56522 (
    .I(net_5),
    .O(net_56522)
  );
  ClkMux inmux_13_31_5_56523 (
    .I(net_5),
    .O(net_56523)
  );
  InMux inmux_13_3_53073_53145 (
    .I(net_53073),
    .O(net_53145)
  );
  InMux inmux_13_3_53074_53142 (
    .I(net_53074),
    .O(net_53142)
  );
  CEMux inmux_13_3_53078_53146 (
    .I(net_53078),
    .O(net_53146)
  );
  InMux inmux_13_3_53092_53143 (
    .I(net_53092),
    .O(net_53143)
  );
  InMux inmux_13_3_53095_53144 (
    .I(net_53095),
    .O(net_53144)
  );
  InMux inmux_13_3_53098_53109 (
    .I(net_53098),
    .O(net_53109)
  );
  ClkMux inmux_13_3_5_53147 (
    .I(net_5),
    .O(net_53147)
  );
  InMux inmux_13_4_53194_53259 (
    .I(net_53194),
    .O(net_53259)
  );
  InMux inmux_13_4_53198_53260 (
    .I(net_53198),
    .O(net_53260)
  );
  InMux inmux_13_4_53198_53265 (
    .I(net_53198),
    .O(net_53265)
  );
  InMux inmux_13_4_53204_53248 (
    .I(net_53204),
    .O(net_53248)
  );
  CEMux inmux_13_4_53208_53269 (
    .I(net_53208),
    .O(net_53269)
  );
  InMux inmux_13_4_53210_53242 (
    .I(net_53210),
    .O(net_53242)
  );
  InMux inmux_13_4_53211_53267 (
    .I(net_53211),
    .O(net_53267)
  );
  InMux inmux_13_4_53213_53255 (
    .I(net_53213),
    .O(net_53255)
  );
  InMux inmux_13_4_53214_53231 (
    .I(net_53214),
    .O(net_53231)
  );
  InMux inmux_13_4_53215_53237 (
    .I(net_53215),
    .O(net_53237)
  );
  InMux inmux_13_4_53221_53225 (
    .I(net_53221),
    .O(net_53225)
  );
  InMux inmux_13_4_53228_53238 (
    .I(net_53228),
    .O(net_53238)
  );
  InMux inmux_13_4_53234_53244 (
    .I(net_53234),
    .O(net_53244)
  );
  InMux inmux_13_4_53240_53250 (
    .I(net_53240),
    .O(net_53250)
  );
  InMux inmux_13_4_53246_53256 (
    .I(net_53246),
    .O(net_53256)
  );
  ClkMux inmux_13_4_5_53270 (
    .I(net_5),
    .O(net_53270)
  );
  InMux inmux_13_8_53682_53722 (
    .I(net_53682),
    .O(net_53722)
  );
  InMux inmux_13_8_53683_53728 (
    .I(net_53683),
    .O(net_53728)
  );
  InMux inmux_13_8_53687_53759 (
    .I(net_53687),
    .O(net_53759)
  );
  InMux inmux_13_8_53688_53741 (
    .I(net_53688),
    .O(net_53741)
  );
  InMux inmux_13_8_53690_53747 (
    .I(net_53690),
    .O(net_53747)
  );
  InMux inmux_13_8_53696_53716 (
    .I(net_53696),
    .O(net_53716)
  );
  InMux inmux_13_8_53712_53735 (
    .I(net_53712),
    .O(net_53735)
  );
  InMux inmux_13_8_53713_53753 (
    .I(net_53713),
    .O(net_53753)
  );
  InMux inmux_13_8_53720_53730 (
    .I(net_53720),
    .O(net_53730)
  );
  InMux inmux_13_8_53726_53736 (
    .I(net_53726),
    .O(net_53736)
  );
  InMux inmux_13_8_53732_53742 (
    .I(net_53732),
    .O(net_53742)
  );
  InMux inmux_13_8_53738_53748 (
    .I(net_53738),
    .O(net_53748)
  );
  InMux inmux_13_8_53744_53754 (
    .I(net_53744),
    .O(net_53754)
  );
  InMux inmux_13_8_53750_53760 (
    .I(net_53750),
    .O(net_53760)
  );
  InMux inmux_13_9_53807_53847 (
    .I(net_53807),
    .O(net_53847)
  );
  InMux inmux_13_9_53809_53876 (
    .I(net_53809),
    .O(net_53876)
  );
  InMux inmux_13_9_53814_53850 (
    .I(net_53814),
    .O(net_53850)
  );
  InMux inmux_13_9_53815_53841 (
    .I(net_53815),
    .O(net_53841)
  );
  InMux inmux_13_9_53815_53846 (
    .I(net_53815),
    .O(net_53846)
  );
  InMux inmux_13_9_53815_53870 (
    .I(net_53815),
    .O(net_53870)
  );
  InMux inmux_13_9_53815_53877 (
    .I(net_53815),
    .O(net_53877)
  );
  InMux inmux_13_9_53817_53853 (
    .I(net_53817),
    .O(net_53853)
  );
  InMux inmux_13_9_53818_53838 (
    .I(net_53818),
    .O(net_53838)
  );
  InMux inmux_13_9_53819_53851 (
    .I(net_53819),
    .O(net_53851)
  );
  InMux inmux_13_9_53820_53871 (
    .I(net_53820),
    .O(net_53871)
  );
  InMux inmux_13_9_53823_53845 (
    .I(net_53823),
    .O(net_53845)
  );
  InMux inmux_13_9_53825_53874 (
    .I(net_53825),
    .O(net_53874)
  );
  InMux inmux_13_9_53827_53852 (
    .I(net_53827),
    .O(net_53852)
  );
  InMux inmux_13_9_53831_53839 (
    .I(net_53831),
    .O(net_53839)
  );
  InMux inmux_13_9_53831_53844 (
    .I(net_53831),
    .O(net_53844)
  );
  InMux inmux_13_9_53831_53868 (
    .I(net_53831),
    .O(net_53868)
  );
  InMux inmux_13_9_53831_53875 (
    .I(net_53831),
    .O(net_53875)
  );
  CEMux inmux_13_9_53832_53884 (
    .I(net_53832),
    .O(net_53884)
  );
  InMux inmux_13_9_53834_53840 (
    .I(net_53834),
    .O(net_53840)
  );
  InMux inmux_13_9_53836_53869 (
    .I(net_53836),
    .O(net_53869)
  );
  ClkMux inmux_13_9_5_53885 (
    .I(net_5),
    .O(net_53885)
  );
  InMux inmux_14_10_57763_57833 (
    .I(net_57763),
    .O(net_57833)
  );
  InMux inmux_14_10_57764_57836 (
    .I(net_57764),
    .O(net_57836)
  );
  InMux inmux_14_10_57776_57834 (
    .I(net_57776),
    .O(net_57834)
  );
  InMux inmux_14_10_57779_57835 (
    .I(net_57779),
    .O(net_57835)
  );
  InMux inmux_14_11_57884_57915 (
    .I(net_57884),
    .O(net_57915)
  );
  InMux inmux_14_11_57885_57940 (
    .I(net_57885),
    .O(net_57940)
  );
  InMux inmux_14_11_57887_57938 (
    .I(net_57887),
    .O(net_57938)
  );
  InMux inmux_14_11_57888_57941 (
    .I(net_57888),
    .O(net_57941)
  );
  InMux inmux_14_11_57888_57944 (
    .I(net_57888),
    .O(net_57944)
  );
  InMux inmux_14_11_57890_57928 (
    .I(net_57890),
    .O(net_57928)
  );
  InMux inmux_14_11_57890_57952 (
    .I(net_57890),
    .O(net_57952)
  );
  InMux inmux_14_11_57893_57929 (
    .I(net_57893),
    .O(net_57929)
  );
  InMux inmux_14_11_57893_57939 (
    .I(net_57893),
    .O(net_57939)
  );
  InMux inmux_14_11_57897_57959 (
    .I(net_57897),
    .O(net_57959)
  );
  InMux inmux_14_11_57899_57926 (
    .I(net_57899),
    .O(net_57926)
  );
  InMux inmux_14_11_57900_57920 (
    .I(net_57900),
    .O(net_57920)
  );
  InMux inmux_14_11_57902_57927 (
    .I(net_57902),
    .O(net_57927)
  );
  InMux inmux_14_11_57903_57933 (
    .I(net_57903),
    .O(net_57933)
  );
  ClkMux inmux_14_11_5_57961 (
    .I(net_5),
    .O(net_57961)
  );
  CEMux inmux_14_11_8_57960 (
    .I(net_8),
    .O(net_57960)
  );
  CEMux inmux_14_12_58006_58083 (
    .I(net_58006),
    .O(net_58083)
  );
  InMux inmux_14_12_58007_58076 (
    .I(net_58007),
    .O(net_58076)
  );
  InMux inmux_14_12_58012_58038 (
    .I(net_58012),
    .O(net_58038)
  );
  InMux inmux_14_12_58012_58052 (
    .I(net_58012),
    .O(net_58052)
  );
  InMux inmux_14_12_58012_58055 (
    .I(net_58012),
    .O(net_58055)
  );
  InMux inmux_14_12_58012_58081 (
    .I(net_58012),
    .O(net_58081)
  );
  InMux inmux_14_12_58013_58082 (
    .I(net_58013),
    .O(net_58082)
  );
  InMux inmux_14_12_58014_58050 (
    .I(net_58014),
    .O(net_58050)
  );
  InMux inmux_14_12_58015_58058 (
    .I(net_58015),
    .O(net_58058)
  );
  InMux inmux_14_12_58018_58043 (
    .I(net_58018),
    .O(net_58043)
  );
  InMux inmux_14_12_58019_58037 (
    .I(net_58019),
    .O(net_58037)
  );
  InMux inmux_14_12_58021_58064 (
    .I(net_58021),
    .O(net_58064)
  );
  InMux inmux_14_12_58023_58040 (
    .I(net_58023),
    .O(net_58040)
  );
  InMux inmux_14_12_58024_58051 (
    .I(net_58024),
    .O(net_58051)
  );
  InMux inmux_14_12_58026_58049 (
    .I(net_58026),
    .O(net_58049)
  );
  InMux inmux_14_12_58026_58056 (
    .I(net_58026),
    .O(net_58056)
  );
  InMux inmux_14_12_58027_58079 (
    .I(net_58027),
    .O(net_58079)
  );
  InMux inmux_14_12_58031_58080 (
    .I(net_58031),
    .O(net_58080)
  );
  InMux inmux_14_12_58034_58057 (
    .I(net_58034),
    .O(net_58057)
  );
  InMux inmux_14_12_58034_58067 (
    .I(net_58034),
    .O(net_58067)
  );
  InMux inmux_14_12_58035_58039 (
    .I(net_58035),
    .O(net_58039)
  );
  ClkMux inmux_14_12_5_58084 (
    .I(net_5),
    .O(net_58084)
  );
  InMux inmux_14_13_58128_58166 (
    .I(net_58128),
    .O(net_58166)
  );
  InMux inmux_14_13_58129_58179 (
    .I(net_58129),
    .O(net_58179)
  );
  InMux inmux_14_13_58130_58178 (
    .I(net_58130),
    .O(net_58178)
  );
  InMux inmux_14_13_58133_58196 (
    .I(net_58133),
    .O(net_58196)
  );
  InMux inmux_14_13_58134_58192 (
    .I(net_58134),
    .O(net_58192)
  );
  InMux inmux_14_13_58135_58173 (
    .I(net_58135),
    .O(net_58173)
  );
  InMux inmux_14_13_58136_58186 (
    .I(net_58136),
    .O(net_58186)
  );
  InMux inmux_14_13_58137_58197 (
    .I(net_58137),
    .O(net_58197)
  );
  InMux inmux_14_13_58138_58181 (
    .I(net_58138),
    .O(net_58181)
  );
  InMux inmux_14_13_58140_58169 (
    .I(net_58140),
    .O(net_58169)
  );
  InMux inmux_14_13_58140_58184 (
    .I(net_58140),
    .O(net_58184)
  );
  InMux inmux_14_13_58140_58193 (
    .I(net_58140),
    .O(net_58193)
  );
  InMux inmux_14_13_58141_58185 (
    .I(net_58141),
    .O(net_58185)
  );
  InMux inmux_14_13_58142_58160 (
    .I(net_58142),
    .O(net_58160)
  );
  InMux inmux_14_13_58144_58168 (
    .I(net_58144),
    .O(net_58168)
  );
  InMux inmux_14_13_58145_58191 (
    .I(net_58145),
    .O(net_58191)
  );
  InMux inmux_14_13_58147_58203 (
    .I(net_58147),
    .O(net_58203)
  );
  InMux inmux_14_13_58148_58187 (
    .I(net_58148),
    .O(net_58187)
  );
  InMux inmux_14_13_58149_58172 (
    .I(net_58149),
    .O(net_58172)
  );
  InMux inmux_14_13_58150_58190 (
    .I(net_58150),
    .O(net_58190)
  );
  InMux inmux_14_13_58151_58199 (
    .I(net_58151),
    .O(net_58199)
  );
  InMux inmux_14_13_58152_58198 (
    .I(net_58152),
    .O(net_58198)
  );
  CEMux inmux_14_13_58154_58206 (
    .I(net_58154),
    .O(net_58206)
  );
  InMux inmux_14_13_58155_58180 (
    .I(net_58155),
    .O(net_58180)
  );
  InMux inmux_14_13_58156_58174 (
    .I(net_58156),
    .O(net_58174)
  );
  InMux inmux_14_13_58157_58175 (
    .I(net_58157),
    .O(net_58175)
  );
  InMux inmux_14_13_58158_58167 (
    .I(net_58158),
    .O(net_58167)
  );
  ClkMux inmux_14_13_5_58207 (
    .I(net_5),
    .O(net_58207)
  );
  InMux inmux_14_14_58258_58286 (
    .I(net_58258),
    .O(net_58286)
  );
  InMux inmux_14_14_58260_58298 (
    .I(net_58260),
    .O(net_58298)
  );
  InMux inmux_14_14_58260_58325 (
    .I(net_58260),
    .O(net_58325)
  );
  InMux inmux_14_14_58261_58295 (
    .I(net_58261),
    .O(net_58295)
  );
  InMux inmux_14_14_58262_58310 (
    .I(net_58262),
    .O(net_58310)
  );
  InMux inmux_14_14_58263_58285 (
    .I(net_58263),
    .O(net_58285)
  );
  InMux inmux_14_14_58264_58327 (
    .I(net_58264),
    .O(net_58327)
  );
  InMux inmux_14_14_58270_58319 (
    .I(net_58270),
    .O(net_58319)
  );
  InMux inmux_14_14_58272_58297 (
    .I(net_58272),
    .O(net_58297)
  );
  InMux inmux_14_14_58273_58284 (
    .I(net_58273),
    .O(net_58284)
  );
  InMux inmux_14_14_58274_58315 (
    .I(net_58274),
    .O(net_58315)
  );
  InMux inmux_14_14_58276_58296 (
    .I(net_58276),
    .O(net_58296)
  );
  InMux inmux_14_14_58277_58283 (
    .I(net_58277),
    .O(net_58283)
  );
  InMux inmux_14_14_58277_58290 (
    .I(net_58277),
    .O(net_58290)
  );
  InMux inmux_14_14_58277_58309 (
    .I(net_58277),
    .O(net_58309)
  );
  InMux inmux_14_14_58279_58302 (
    .I(net_58279),
    .O(net_58302)
  );
  InMux inmux_14_14_58279_58328 (
    .I(net_58279),
    .O(net_58328)
  );
  InMux inmux_14_14_58280_58291 (
    .I(net_58280),
    .O(net_58291)
  );
  InMux inmux_14_14_58281_58326 (
    .I(net_58281),
    .O(net_58326)
  );
  ClkMux inmux_14_14_5_58330 (
    .I(net_5),
    .O(net_58330)
  );
  CEMux inmux_14_14_8_58329 (
    .I(net_8),
    .O(net_58329)
  );
  InMux inmux_14_15_58382_58427 (
    .I(net_58382),
    .O(net_58427)
  );
  InMux inmux_14_15_58383_58414 (
    .I(net_58383),
    .O(net_58414)
  );
  InMux inmux_14_15_58383_58438 (
    .I(net_58383),
    .O(net_58438)
  );
  InMux inmux_14_15_58386_58425 (
    .I(net_58386),
    .O(net_58425)
  );
  InMux inmux_14_15_58387_58426 (
    .I(net_58387),
    .O(net_58426)
  );
  CEMux inmux_14_15_58391_58452 (
    .I(net_58391),
    .O(net_58452)
  );
  InMux inmux_14_15_58392_58407 (
    .I(net_58392),
    .O(net_58407)
  );
  InMux inmux_14_15_58395_58420 (
    .I(net_58395),
    .O(net_58420)
  );
  InMux inmux_14_15_58396_58448 (
    .I(net_58396),
    .O(net_58448)
  );
  InMux inmux_14_15_58397_58424 (
    .I(net_58397),
    .O(net_58424)
  );
  InMux inmux_14_15_58398_58415 (
    .I(net_58398),
    .O(net_58415)
  );
  InMux inmux_14_15_58402_58432 (
    .I(net_58402),
    .O(net_58432)
  );
  InMux inmux_14_15_58403_58445 (
    .I(net_58403),
    .O(net_58445)
  );
  InMux inmux_14_15_58404_58437 (
    .I(net_58404),
    .O(net_58437)
  );
  ClkMux inmux_14_15_5_58453 (
    .I(net_5),
    .O(net_58453)
  );
  CEMux inmux_14_16_58498_58575 (
    .I(net_58498),
    .O(net_58575)
  );
  InMux inmux_14_16_58500_58550 (
    .I(net_58500),
    .O(net_58550)
  );
  InMux inmux_14_16_58501_58568 (
    .I(net_58501),
    .O(net_58568)
  );
  InMux inmux_14_16_58504_58571 (
    .I(net_58504),
    .O(net_58571)
  );
  InMux inmux_14_16_58509_58538 (
    .I(net_58509),
    .O(net_58538)
  );
  InMux inmux_14_16_58511_58531 (
    .I(net_58511),
    .O(net_58531)
  );
  InMux inmux_14_16_58513_58559 (
    .I(net_58513),
    .O(net_58559)
  );
  InMux inmux_14_16_58517_58537 (
    .I(net_58517),
    .O(net_58537)
  );
  InMux inmux_14_16_58518_58555 (
    .I(net_58518),
    .O(net_58555)
  );
  InMux inmux_14_16_58520_58535 (
    .I(net_58520),
    .O(net_58535)
  );
  InMux inmux_14_16_58521_58536 (
    .I(net_58521),
    .O(net_58536)
  );
  InMux inmux_14_16_58523_58553 (
    .I(net_58523),
    .O(net_58553)
  );
  ClkMux inmux_14_16_5_58576 (
    .I(net_5),
    .O(net_58576)
  );
  InMux inmux_14_17_58620_58658 (
    .I(net_58620),
    .O(net_58658)
  );
  CEMux inmux_14_17_58630_58698 (
    .I(net_58630),
    .O(net_58698)
  );
  InMux inmux_14_17_58633_58682 (
    .I(net_58633),
    .O(net_58682)
  );
  InMux inmux_14_17_58644_58671 (
    .I(net_58644),
    .O(net_58671)
  );
  InMux inmux_14_17_58644_58685 (
    .I(net_58644),
    .O(net_58685)
  );
  InMux inmux_14_17_58645_58665 (
    .I(net_58645),
    .O(net_58665)
  );
  InMux inmux_14_17_58650_58695 (
    .I(net_58650),
    .O(net_58695)
  );
  ClkMux inmux_14_17_5_58699 (
    .I(net_5),
    .O(net_58699)
  );
  InMux inmux_14_18_58745_58817 (
    .I(net_58745),
    .O(net_58817)
  );
  InMux inmux_14_18_58747_58800 (
    .I(net_58747),
    .O(net_58800)
  );
  InMux inmux_14_18_58749_58781 (
    .I(net_58749),
    .O(net_58781)
  );
  InMux inmux_14_18_58753_58820 (
    .I(net_58753),
    .O(net_58820)
  );
  InMux inmux_14_18_58758_58808 (
    .I(net_58758),
    .O(net_58808)
  );
  InMux inmux_14_18_58759_58819 (
    .I(net_58759),
    .O(net_58819)
  );
  InMux inmux_14_18_58760_58799 (
    .I(net_58760),
    .O(net_58799)
  );
  InMux inmux_14_18_58760_58818 (
    .I(net_58760),
    .O(net_58818)
  );
  InMux inmux_14_18_58761_58776 (
    .I(net_58761),
    .O(net_58776)
  );
  InMux inmux_14_18_58761_58793 (
    .I(net_58761),
    .O(net_58793)
  );
  InMux inmux_14_18_58763_58778 (
    .I(net_58763),
    .O(net_58778)
  );
  InMux inmux_14_18_58764_58801 (
    .I(net_58764),
    .O(net_58801)
  );
  InMux inmux_14_18_58766_58802 (
    .I(net_58766),
    .O(net_58802)
  );
  InMux inmux_14_18_58767_58796 (
    .I(net_58767),
    .O(net_58796)
  );
  CEMux inmux_14_18_58769_58821 (
    .I(net_58769),
    .O(net_58821)
  );
  ClkMux inmux_14_18_5_58822 (
    .I(net_5),
    .O(net_58822)
  );
  InMux inmux_14_19_58865_58941 (
    .I(net_58865),
    .O(net_58941)
  );
  InMux inmux_14_19_58867_58907 (
    .I(net_58867),
    .O(net_58907)
  );
  InMux inmux_14_19_58873_58906 (
    .I(net_58873),
    .O(net_58906)
  );
  InMux inmux_14_19_58875_58899 (
    .I(net_58875),
    .O(net_58899)
  );
  InMux inmux_14_19_58877_58935 (
    .I(net_58877),
    .O(net_58935)
  );
  InMux inmux_14_19_58884_58904 (
    .I(net_58884),
    .O(net_58904)
  );
  InMux inmux_14_19_58892_58936 (
    .I(net_58892),
    .O(net_58936)
  );
  InMux inmux_14_19_58892_58943 (
    .I(net_58892),
    .O(net_58943)
  );
  InMux inmux_14_19_58894_58905 (
    .I(net_58894),
    .O(net_58905)
  );
  ClkMux inmux_14_19_5_58945 (
    .I(net_5),
    .O(net_58945)
  );
  CEMux inmux_14_19_6_58944 (
    .I(net_6),
    .O(net_58944)
  );
  InMux inmux_14_20_58988_59035 (
    .I(net_58988),
    .O(net_59035)
  );
  InMux inmux_14_20_58990_59054 (
    .I(net_58990),
    .O(net_59054)
  );
  InMux inmux_14_20_58991_59027 (
    .I(net_58991),
    .O(net_59027)
  );
  InMux inmux_14_20_58992_59066 (
    .I(net_58992),
    .O(net_59066)
  );
  InMux inmux_14_20_58993_59046 (
    .I(net_58993),
    .O(net_59046)
  );
  InMux inmux_14_20_58994_59052 (
    .I(net_58994),
    .O(net_59052)
  );
  InMux inmux_14_20_58995_59063 (
    .I(net_58995),
    .O(net_59063)
  );
  CEMux inmux_14_20_58999_59067 (
    .I(net_58999),
    .O(net_59067)
  );
  InMux inmux_14_20_59002_59053 (
    .I(net_59002),
    .O(net_59053)
  );
  InMux inmux_14_20_59004_59064 (
    .I(net_59004),
    .O(net_59064)
  );
  InMux inmux_14_20_59005_59051 (
    .I(net_59005),
    .O(net_59051)
  );
  InMux inmux_14_20_59014_59029 (
    .I(net_59014),
    .O(net_59029)
  );
  InMux inmux_14_20_59016_59065 (
    .I(net_59016),
    .O(net_59065)
  );
  InMux inmux_14_20_59017_59023 (
    .I(net_59017),
    .O(net_59023)
  );
  ClkMux inmux_14_20_5_59068 (
    .I(net_5),
    .O(net_59068)
  );
  InMux inmux_14_21_59140_59187 (
    .I(net_59140),
    .O(net_59187)
  );
  ClkMux inmux_14_21_5_59191 (
    .I(net_5),
    .O(net_59191)
  );
  CEMux inmux_14_21_6_59190 (
    .I(net_6),
    .O(net_59190)
  );
  InMux inmux_14_26_59735_59778 (
    .I(net_59735),
    .O(net_59778)
  );
  InMux inmux_14_26_59735_59783 (
    .I(net_59735),
    .O(net_59783)
  );
  CEMux inmux_14_26_59737_59805 (
    .I(net_59737),
    .O(net_59805)
  );
  InMux inmux_14_26_59753_59785 (
    .I(net_59753),
    .O(net_59785)
  );
  ClkMux inmux_14_26_5_59806 (
    .I(net_5),
    .O(net_59806)
  );
  InMux inmux_14_27_59851_59913 (
    .I(net_59851),
    .O(net_59913)
  );
  InMux inmux_14_27_59851_59915 (
    .I(net_59851),
    .O(net_59915)
  );
  InMux inmux_14_27_59859_59914 (
    .I(net_59859),
    .O(net_59914)
  );
  InMux inmux_14_27_59862_59891 (
    .I(net_59862),
    .O(net_59891)
  );
  CEMux inmux_14_27_59867_59928 (
    .I(net_59867),
    .O(net_59928)
  );
  InMux inmux_14_27_59869_59889 (
    .I(net_59869),
    .O(net_59889)
  );
  InMux inmux_14_27_59870_59888 (
    .I(net_59870),
    .O(net_59888)
  );
  InMux inmux_14_27_59875_59895 (
    .I(net_59875),
    .O(net_59895)
  );
  InMux inmux_14_27_59879_59890 (
    .I(net_59879),
    .O(net_59890)
  );
  ClkMux inmux_14_27_5_59929 (
    .I(net_5),
    .O(net_59929)
  );
  InMux inmux_14_28_59984_60011 (
    .I(net_59984),
    .O(net_60011)
  );
  InMux inmux_14_28_59988_60014 (
    .I(net_59988),
    .O(net_60014)
  );
  InMux inmux_14_2_56776_56840 (
    .I(net_56776),
    .O(net_56840)
  );
  InMux inmux_14_2_56776_56843 (
    .I(net_56776),
    .O(net_56843)
  );
  InMux inmux_14_2_56777_56839 (
    .I(net_56777),
    .O(net_56839)
  );
  InMux inmux_14_2_56780_56845 (
    .I(net_56780),
    .O(net_56845)
  );
  InMux inmux_14_2_56785_56838 (
    .I(net_56785),
    .O(net_56838)
  );
  InMux inmux_14_2_56790_56821 (
    .I(net_56790),
    .O(net_56821)
  );
  InMux inmux_14_2_56790_56828 (
    .I(net_56790),
    .O(net_56828)
  );
  InMux inmux_14_2_56793_56825 (
    .I(net_56793),
    .O(net_56825)
  );
  InMux inmux_14_2_56793_56844 (
    .I(net_56793),
    .O(net_56844)
  );
  InMux inmux_14_2_56800_56827 (
    .I(net_56800),
    .O(net_56827)
  );
  InMux inmux_14_2_56800_56846 (
    .I(net_56800),
    .O(net_56846)
  );
  InMux inmux_14_2_56805_56819 (
    .I(net_56805),
    .O(net_56819)
  );
  InMux inmux_14_2_56805_56826 (
    .I(net_56805),
    .O(net_56826)
  );
  InMux inmux_14_3_56897_56942 (
    .I(net_56897),
    .O(net_56942)
  );
  InMux inmux_14_3_56897_56949 (
    .I(net_56897),
    .O(net_56949)
  );
  InMux inmux_14_3_56898_56955 (
    .I(net_56898),
    .O(net_56955)
  );
  InMux inmux_14_3_56899_56956 (
    .I(net_56899),
    .O(net_56956)
  );
  InMux inmux_14_3_56904_56943 (
    .I(net_56904),
    .O(net_56943)
  );
  InMux inmux_14_3_56904_56972 (
    .I(net_56904),
    .O(net_56972)
  );
  InMux inmux_14_3_56905_56931 (
    .I(net_56905),
    .O(net_56931)
  );
  InMux inmux_14_3_56905_56962 (
    .I(net_56905),
    .O(net_56962)
  );
  InMux inmux_14_3_56905_56967 (
    .I(net_56905),
    .O(net_56967)
  );
  InMux inmux_14_3_56906_56951 (
    .I(net_56906),
    .O(net_56951)
  );
  InMux inmux_14_3_56908_56961 (
    .I(net_56908),
    .O(net_56961)
  );
  InMux inmux_14_3_56909_56950 (
    .I(net_56909),
    .O(net_56950)
  );
  InMux inmux_14_3_56911_56960 (
    .I(net_56911),
    .O(net_56960)
  );
  InMux inmux_14_3_56912_56954 (
    .I(net_56912),
    .O(net_56954)
  );
  InMux inmux_14_3_56914_56948 (
    .I(net_56914),
    .O(net_56948)
  );
  InMux inmux_14_3_56915_56932 (
    .I(net_56915),
    .O(net_56932)
  );
  InMux inmux_14_3_56915_56968 (
    .I(net_56915),
    .O(net_56968)
  );
  InMux inmux_14_3_56916_56933 (
    .I(net_56916),
    .O(net_56933)
  );
  InMux inmux_14_3_56916_56969 (
    .I(net_56916),
    .O(net_56969)
  );
  InMux inmux_14_3_56917_56937 (
    .I(net_56917),
    .O(net_56937)
  );
  InMux inmux_14_3_56917_56939 (
    .I(net_56917),
    .O(net_56939)
  );
  InMux inmux_14_3_56920_56938 (
    .I(net_56920),
    .O(net_56938)
  );
  InMux inmux_14_3_56921_56957 (
    .I(net_56921),
    .O(net_56957)
  );
  CEMux inmux_14_3_56924_56976 (
    .I(net_56924),
    .O(net_56976)
  );
  InMux inmux_14_3_56928_56930 (
    .I(net_56928),
    .O(net_56930)
  );
  InMux inmux_14_3_56928_56963 (
    .I(net_56928),
    .O(net_56963)
  );
  InMux inmux_14_3_56928_56966 (
    .I(net_56928),
    .O(net_56966)
  );
  ClkMux inmux_14_3_5_56977 (
    .I(net_5),
    .O(net_56977)
  );
  InMux inmux_14_4_57023_57078 (
    .I(net_57023),
    .O(net_57078)
  );
  InMux inmux_14_4_57027_57083 (
    .I(net_57027),
    .O(net_57083)
  );
  InMux inmux_14_4_57028_57056 (
    .I(net_57028),
    .O(net_57056)
  );
  InMux inmux_14_4_57028_57059 (
    .I(net_57028),
    .O(net_57059)
  );
  InMux inmux_14_4_57028_57080 (
    .I(net_57028),
    .O(net_57080)
  );
  InMux inmux_14_4_57028_57097 (
    .I(net_57028),
    .O(net_57097)
  );
  InMux inmux_14_4_57030_57061 (
    .I(net_57030),
    .O(net_57061)
  );
  InMux inmux_14_4_57034_57066 (
    .I(net_57034),
    .O(net_57066)
  );
  CEMux inmux_14_4_57038_57099 (
    .I(net_57038),
    .O(net_57099)
  );
  InMux inmux_14_4_57041_57085 (
    .I(net_57041),
    .O(net_57085)
  );
  InMux inmux_14_4_57044_57054 (
    .I(net_57044),
    .O(net_57054)
  );
  InMux inmux_14_4_57046_57068 (
    .I(net_57046),
    .O(net_57068)
  );
  InMux inmux_14_4_57049_57098 (
    .I(net_57049),
    .O(net_57098)
  );
  InMux inmux_14_4_57051_57053 (
    .I(net_57051),
    .O(net_57053)
  );
  ClkMux inmux_14_4_5_57100 (
    .I(net_5),
    .O(net_57100)
  );
  CEMux inmux_14_7_57391_57468 (
    .I(net_57391),
    .O(net_57468)
  );
  InMux inmux_14_7_57403_57428 (
    .I(net_57403),
    .O(net_57428)
  );
  InMux inmux_14_7_57403_57464 (
    .I(net_57403),
    .O(net_57464)
  );
  InMux inmux_14_7_57410_57461 (
    .I(net_57410),
    .O(net_57461)
  );
  InMux inmux_14_7_57412_57459 (
    .I(net_57412),
    .O(net_57459)
  );
  InMux inmux_14_7_57414_57458 (
    .I(net_57414),
    .O(net_57458)
  );
  InMux inmux_14_7_57415_57430 (
    .I(net_57415),
    .O(net_57430)
  );
  InMux inmux_14_7_57415_57466 (
    .I(net_57415),
    .O(net_57466)
  );
  InMux inmux_14_7_57418_57460 (
    .I(net_57418),
    .O(net_57460)
  );
  ClkMux inmux_14_7_5_57469 (
    .I(net_5),
    .O(net_57469)
  );
  InMux inmux_14_8_57515_57584 (
    .I(net_57515),
    .O(net_57584)
  );
  InMux inmux_14_8_57518_57588 (
    .I(net_57518),
    .O(net_57588)
  );
  InMux inmux_14_8_57523_57581 (
    .I(net_57523),
    .O(net_57581)
  );
  InMux inmux_14_8_57526_57572 (
    .I(net_57526),
    .O(net_57572)
  );
  InMux inmux_14_8_57526_57575 (
    .I(net_57526),
    .O(net_57575)
  );
  InMux inmux_14_8_57527_57571 (
    .I(net_57527),
    .O(net_57571)
  );
  InMux inmux_14_8_57528_57578 (
    .I(net_57528),
    .O(net_57578)
  );
  InMux inmux_14_8_57528_57583 (
    .I(net_57528),
    .O(net_57583)
  );
  InMux inmux_14_8_57528_57590 (
    .I(net_57528),
    .O(net_57590)
  );
  InMux inmux_14_8_57529_57589 (
    .I(net_57529),
    .O(net_57589)
  );
  InMux inmux_14_8_57535_57582 (
    .I(net_57535),
    .O(net_57582)
  );
  InMux inmux_14_8_57535_57587 (
    .I(net_57535),
    .O(net_57587)
  );
  InMux inmux_14_8_57536_57570 (
    .I(net_57536),
    .O(net_57570)
  );
  CEMux inmux_14_8_57539_57591 (
    .I(net_57539),
    .O(net_57591)
  );
  InMux inmux_14_8_57541_57569 (
    .I(net_57541),
    .O(net_57569)
  );
  InMux inmux_14_8_57543_57576 (
    .I(net_57543),
    .O(net_57576)
  );
  ClkMux inmux_14_8_5_57592 (
    .I(net_5),
    .O(net_57592)
  );
  InMux inmux_14_9_57635_57699 (
    .I(net_57635),
    .O(net_57699)
  );
  InMux inmux_14_9_57636_57681 (
    .I(net_57636),
    .O(net_57681)
  );
  InMux inmux_14_9_57640_57710 (
    .I(net_57640),
    .O(net_57710)
  );
  InMux inmux_14_9_57641_57694 (
    .I(net_57641),
    .O(net_57694)
  );
  InMux inmux_14_9_57642_57705 (
    .I(net_57642),
    .O(net_57705)
  );
  InMux inmux_14_9_57643_57676 (
    .I(net_57643),
    .O(net_57676)
  );
  InMux inmux_14_9_57647_57669 (
    .I(net_57647),
    .O(net_57669)
  );
  InMux inmux_14_9_57649_57688 (
    .I(net_57649),
    .O(net_57688)
  );
  InMux inmux_14_9_57652_57693 (
    .I(net_57652),
    .O(net_57693)
  );
  InMux inmux_14_9_57652_57700 (
    .I(net_57652),
    .O(net_57700)
  );
  InMux inmux_14_9_57652_57712 (
    .I(net_57652),
    .O(net_57712)
  );
  InMux inmux_14_9_57660_57675 (
    .I(net_57660),
    .O(net_57675)
  );
  InMux inmux_14_9_57660_57682 (
    .I(net_57660),
    .O(net_57682)
  );
  InMux inmux_14_9_57660_57687 (
    .I(net_57660),
    .O(net_57687)
  );
  InMux inmux_14_9_57660_57706 (
    .I(net_57660),
    .O(net_57706)
  );
  InMux inmux_14_9_57673_57683 (
    .I(net_57673),
    .O(net_57683)
  );
  InMux inmux_14_9_57679_57689 (
    .I(net_57679),
    .O(net_57689)
  );
  InMux inmux_14_9_57685_57695 (
    .I(net_57685),
    .O(net_57695)
  );
  InMux inmux_14_9_57691_57701 (
    .I(net_57691),
    .O(net_57701)
  );
  InMux inmux_14_9_57697_57707 (
    .I(net_57697),
    .O(net_57707)
  );
  InMux inmux_14_9_57703_57713 (
    .I(net_57703),
    .O(net_57713)
  );
  ClkMux inmux_15_10_5_61668 (
    .I(net_5),
    .O(net_61668)
  );
  InMux inmux_15_10_61588_61623 (
    .I(net_61588),
    .O(net_61623)
  );
  InMux inmux_15_10_61591_61651 (
    .I(net_61591),
    .O(net_61651)
  );
  InMux inmux_15_10_61592_61654 (
    .I(net_61592),
    .O(net_61654)
  );
  InMux inmux_15_10_61594_61657 (
    .I(net_61594),
    .O(net_61657)
  );
  InMux inmux_15_10_61596_61653 (
    .I(net_61596),
    .O(net_61653)
  );
  InMux inmux_15_10_61598_61634 (
    .I(net_61598),
    .O(net_61634)
  );
  CEMux inmux_15_10_61599_61667 (
    .I(net_61599),
    .O(net_61667)
  );
  InMux inmux_15_10_61600_61648 (
    .I(net_61600),
    .O(net_61648)
  );
  InMux inmux_15_10_61601_61645 (
    .I(net_61601),
    .O(net_61645)
  );
  InMux inmux_15_10_61602_61629 (
    .I(net_61602),
    .O(net_61629)
  );
  InMux inmux_15_10_61609_61658 (
    .I(net_61609),
    .O(net_61658)
  );
  InMux inmux_15_10_61610_61647 (
    .I(net_61610),
    .O(net_61647)
  );
  InMux inmux_15_10_61613_61652 (
    .I(net_61613),
    .O(net_61652)
  );
  InMux inmux_15_10_61616_61646 (
    .I(net_61616),
    .O(net_61646)
  );
  InMux inmux_15_10_61617_61659 (
    .I(net_61617),
    .O(net_61659)
  );
  InMux inmux_15_10_61626_61636 (
    .I(net_61626),
    .O(net_61636)
  );
  ClkMux inmux_15_11_5_61791 (
    .I(net_5),
    .O(net_61791)
  );
  InMux inmux_15_11_61715_61770 (
    .I(net_61715),
    .O(net_61770)
  );
  InMux inmux_15_11_61716_61752 (
    .I(net_61716),
    .O(net_61752)
  );
  InMux inmux_15_11_61717_61782 (
    .I(net_61717),
    .O(net_61782)
  );
  InMux inmux_15_11_61719_61769 (
    .I(net_61719),
    .O(net_61769)
  );
  InMux inmux_15_11_61724_61746 (
    .I(net_61724),
    .O(net_61746)
  );
  InMux inmux_15_11_61726_61775 (
    .I(net_61726),
    .O(net_61775)
  );
  InMux inmux_15_11_61728_61776 (
    .I(net_61728),
    .O(net_61776)
  );
  CEMux inmux_15_11_61729_61790 (
    .I(net_61729),
    .O(net_61790)
  );
  InMux inmux_15_11_61730_61781 (
    .I(net_61730),
    .O(net_61781)
  );
  InMux inmux_15_11_61731_61758 (
    .I(net_61731),
    .O(net_61758)
  );
  InMux inmux_15_11_61735_61788 (
    .I(net_61735),
    .O(net_61788)
  );
  InMux inmux_15_11_61736_61763 (
    .I(net_61736),
    .O(net_61763)
  );
  InMux inmux_15_11_61737_61764 (
    .I(net_61737),
    .O(net_61764)
  );
  InMux inmux_15_11_61738_61787 (
    .I(net_61738),
    .O(net_61787)
  );
  InMux inmux_15_11_61739_61745 (
    .I(net_61739),
    .O(net_61745)
  );
  InMux inmux_15_11_61740_61751 (
    .I(net_61740),
    .O(net_61751)
  );
  InMux inmux_15_11_61741_61757 (
    .I(net_61741),
    .O(net_61757)
  );
  InMux inmux_15_11_61743_61753 (
    .I(net_61743),
    .O(net_61753)
  );
  InMux inmux_15_11_61749_61759 (
    .I(net_61749),
    .O(net_61759)
  );
  InMux inmux_15_11_61755_61765 (
    .I(net_61755),
    .O(net_61765)
  );
  InMux inmux_15_11_61761_61771 (
    .I(net_61761),
    .O(net_61771)
  );
  InMux inmux_15_11_61767_61777 (
    .I(net_61767),
    .O(net_61777)
  );
  InMux inmux_15_11_61773_61783 (
    .I(net_61773),
    .O(net_61783)
  );
  InMux inmux_15_11_61779_61789 (
    .I(net_61779),
    .O(net_61789)
  );
  ClkMux inmux_15_12_5_61914 (
    .I(net_5),
    .O(net_61914)
  );
  InMux inmux_15_12_61829_61870 (
    .I(net_61829),
    .O(net_61870)
  );
  InMux inmux_15_12_61837_61880 (
    .I(net_61837),
    .O(net_61880)
  );
  InMux inmux_15_12_61838_61874 (
    .I(net_61838),
    .O(net_61874)
  );
  InMux inmux_15_12_61841_61904 (
    .I(net_61841),
    .O(net_61904)
  );
  InMux inmux_15_12_61842_61892 (
    .I(net_61842),
    .O(net_61892)
  );
  CEMux inmux_15_12_61845_61913 (
    .I(net_61845),
    .O(net_61913)
  );
  InMux inmux_15_12_61850_61881 (
    .I(net_61850),
    .O(net_61881)
  );
  InMux inmux_15_12_61851_61875 (
    .I(net_61851),
    .O(net_61875)
  );
  InMux inmux_15_12_61852_61886 (
    .I(net_61852),
    .O(net_61886)
  );
  InMux inmux_15_12_61854_61869 (
    .I(net_61854),
    .O(net_61869)
  );
  InMux inmux_15_12_61855_61909 (
    .I(net_61855),
    .O(net_61909)
  );
  InMux inmux_15_12_61856_61893 (
    .I(net_61856),
    .O(net_61893)
  );
  InMux inmux_15_12_61857_61887 (
    .I(net_61857),
    .O(net_61887)
  );
  InMux inmux_15_12_61860_61868 (
    .I(net_61860),
    .O(net_61868)
  );
  InMux inmux_15_12_61861_61898 (
    .I(net_61861),
    .O(net_61898)
  );
  InMux inmux_15_12_61862_61899 (
    .I(net_61862),
    .O(net_61899)
  );
  InMux inmux_15_12_61863_61905 (
    .I(net_61863),
    .O(net_61905)
  );
  InMux inmux_15_12_61864_61911 (
    .I(net_61864),
    .O(net_61911)
  );
  InMux inmux_15_12_61866_61876 (
    .I(net_61866),
    .O(net_61876)
  );
  InMux inmux_15_12_61872_61882 (
    .I(net_61872),
    .O(net_61882)
  );
  InMux inmux_15_12_61878_61888 (
    .I(net_61878),
    .O(net_61888)
  );
  InMux inmux_15_12_61884_61894 (
    .I(net_61884),
    .O(net_61894)
  );
  InMux inmux_15_12_61890_61900 (
    .I(net_61890),
    .O(net_61900)
  );
  InMux inmux_15_12_61896_61906 (
    .I(net_61896),
    .O(net_61906)
  );
  InMux inmux_15_12_61902_61912 (
    .I(net_61902),
    .O(net_61912)
  );
  InMux inmux_15_13_61957_62028 (
    .I(net_61957),
    .O(net_62028)
  );
  InMux inmux_15_13_61961_61992 (
    .I(net_61961),
    .O(net_61992)
  );
  InMux inmux_15_13_61962_62017 (
    .I(net_61962),
    .O(net_62017)
  );
  InMux inmux_15_13_61963_61997 (
    .I(net_61963),
    .O(net_61997)
  );
  InMux inmux_15_13_61965_62010 (
    .I(net_61965),
    .O(net_62010)
  );
  InMux inmux_15_13_61966_61990 (
    .I(net_61966),
    .O(net_61990)
  );
  InMux inmux_15_13_61967_61998 (
    .I(net_61967),
    .O(net_61998)
  );
  InMux inmux_15_13_61968_62021 (
    .I(net_61968),
    .O(net_62021)
  );
  InMux inmux_15_13_61969_61991 (
    .I(net_61969),
    .O(net_61991)
  );
  InMux inmux_15_13_61969_61996 (
    .I(net_61969),
    .O(net_61996)
  );
  InMux inmux_15_13_61969_62005 (
    .I(net_61969),
    .O(net_62005)
  );
  InMux inmux_15_13_61969_62022 (
    .I(net_61969),
    .O(net_62022)
  );
  InMux inmux_15_13_61969_62029 (
    .I(net_61969),
    .O(net_62029)
  );
  InMux inmux_15_13_61970_62002 (
    .I(net_61970),
    .O(net_62002)
  );
  InMux inmux_15_13_61972_62023 (
    .I(net_61972),
    .O(net_62023)
  );
  InMux inmux_15_13_61973_61999 (
    .I(net_61973),
    .O(net_61999)
  );
  InMux inmux_15_13_61974_62003 (
    .I(net_61974),
    .O(net_62003)
  );
  InMux inmux_15_13_61976_61993 (
    .I(net_61976),
    .O(net_61993)
  );
  InMux inmux_15_13_61977_62026 (
    .I(net_61977),
    .O(net_62026)
  );
  InMux inmux_15_13_61978_62027 (
    .I(net_61978),
    .O(net_62027)
  );
  InMux inmux_15_13_61983_62034 (
    .I(net_61983),
    .O(net_62034)
  );
  InMux inmux_15_13_61984_62004 (
    .I(net_61984),
    .O(net_62004)
  );
  InMux inmux_15_13_61985_62020 (
    .I(net_61985),
    .O(net_62020)
  );
  InMux inmux_15_13_61986_62033 (
    .I(net_61986),
    .O(net_62033)
  );
  ClkMux inmux_15_14_5_62160 (
    .I(net_5),
    .O(net_62160)
  );
  InMux inmux_15_14_62081_62145 (
    .I(net_62081),
    .O(net_62145)
  );
  InMux inmux_15_14_62082_62139 (
    .I(net_62082),
    .O(net_62139)
  );
  InMux inmux_15_14_62083_62116 (
    .I(net_62083),
    .O(net_62116)
  );
  InMux inmux_15_14_62086_62149 (
    .I(net_62086),
    .O(net_62149)
  );
  InMux inmux_15_14_62089_62132 (
    .I(net_62089),
    .O(net_62132)
  );
  InMux inmux_15_14_62090_62121 (
    .I(net_62090),
    .O(net_62121)
  );
  InMux inmux_15_14_62090_62140 (
    .I(net_62090),
    .O(net_62140)
  );
  InMux inmux_15_14_62090_62155 (
    .I(net_62090),
    .O(net_62155)
  );
  InMux inmux_15_14_62092_62119 (
    .I(net_62092),
    .O(net_62119)
  );
  InMux inmux_15_14_62094_62138 (
    .I(net_62094),
    .O(net_62138)
  );
  InMux inmux_15_14_62095_62125 (
    .I(net_62095),
    .O(net_62125)
  );
  InMux inmux_15_14_62096_62122 (
    .I(net_62096),
    .O(net_62122)
  );
  InMux inmux_15_14_62098_62158 (
    .I(net_62098),
    .O(net_62158)
  );
  InMux inmux_15_14_62100_62137 (
    .I(net_62100),
    .O(net_62137)
  );
  InMux inmux_15_14_62101_62157 (
    .I(net_62101),
    .O(net_62157)
  );
  InMux inmux_15_14_62105_62120 (
    .I(net_62105),
    .O(net_62120)
  );
  InMux inmux_15_14_62111_62156 (
    .I(net_62111),
    .O(net_62156)
  );
  CEMux inmux_15_14_8_62159 (
    .I(net_8),
    .O(net_62159)
  );
  ClkMux inmux_15_15_5_62283 (
    .I(net_5),
    .O(net_62283)
  );
  InMux inmux_15_15_62204_62249 (
    .I(net_62204),
    .O(net_62249)
  );
  InMux inmux_15_15_62206_62268 (
    .I(net_62206),
    .O(net_62268)
  );
  InMux inmux_15_15_62208_62251 (
    .I(net_62208),
    .O(net_62251)
  );
  InMux inmux_15_15_62209_62260 (
    .I(net_62209),
    .O(net_62260)
  );
  InMux inmux_15_15_62210_62280 (
    .I(net_62210),
    .O(net_62280)
  );
  InMux inmux_15_15_62217_62239 (
    .I(net_62217),
    .O(net_62239)
  );
  InMux inmux_15_15_62218_62250 (
    .I(net_62218),
    .O(net_62250)
  );
  InMux inmux_15_15_62220_62263 (
    .I(net_62220),
    .O(net_62263)
  );
  InMux inmux_15_15_62221_62248 (
    .I(net_62221),
    .O(net_62248)
  );
  InMux inmux_15_15_62224_62266 (
    .I(net_62224),
    .O(net_62266)
  );
  InMux inmux_15_15_62227_62256 (
    .I(net_62227),
    .O(net_62256)
  );
  InMux inmux_15_15_62227_62261 (
    .I(net_62227),
    .O(net_62261)
  );
  InMux inmux_15_15_62229_62275 (
    .I(net_62229),
    .O(net_62275)
  );
  InMux inmux_15_15_62230_62243 (
    .I(net_62230),
    .O(net_62243)
  );
  InMux inmux_15_15_62232_62262 (
    .I(net_62232),
    .O(net_62262)
  );
  CEMux inmux_15_15_8_62282 (
    .I(net_8),
    .O(net_62282)
  );
  ClkMux inmux_15_16_5_62406 (
    .I(net_5),
    .O(net_62406)
  );
  InMux inmux_15_16_62327_62377 (
    .I(net_62327),
    .O(net_62377)
  );
  InMux inmux_15_16_62331_62384 (
    .I(net_62331),
    .O(net_62384)
  );
  InMux inmux_15_16_62334_62386 (
    .I(net_62334),
    .O(net_62386)
  );
  CEMux inmux_15_16_62337_62405 (
    .I(net_62337),
    .O(net_62405)
  );
  InMux inmux_15_16_62339_62395 (
    .I(net_62339),
    .O(net_62395)
  );
  InMux inmux_15_16_62340_62396 (
    .I(net_62340),
    .O(net_62396)
  );
  InMux inmux_15_16_62344_62392 (
    .I(net_62344),
    .O(net_62392)
  );
  InMux inmux_15_16_62346_62385 (
    .I(net_62346),
    .O(net_62385)
  );
  InMux inmux_15_16_62348_62383 (
    .I(net_62348),
    .O(net_62383)
  );
  InMux inmux_15_16_62350_62398 (
    .I(net_62350),
    .O(net_62398)
  );
  InMux inmux_15_16_62353_62359 (
    .I(net_62353),
    .O(net_62359)
  );
  InMux inmux_15_16_62353_62378 (
    .I(net_62353),
    .O(net_62378)
  );
  InMux inmux_15_16_62353_62402 (
    .I(net_62353),
    .O(net_62402)
  );
  InMux inmux_15_16_62354_62403 (
    .I(net_62354),
    .O(net_62403)
  );
  InMux inmux_15_16_62356_62360 (
    .I(net_62356),
    .O(net_62360)
  );
  ClkMux inmux_15_17_5_62529 (
    .I(net_5),
    .O(net_62529)
  );
  InMux inmux_15_17_62456_62526 (
    .I(net_62456),
    .O(net_62526)
  );
  InMux inmux_15_17_62457_62502 (
    .I(net_62457),
    .O(net_62502)
  );
  InMux inmux_15_17_62457_62519 (
    .I(net_62457),
    .O(net_62519)
  );
  InMux inmux_15_17_62458_62491 (
    .I(net_62458),
    .O(net_62491)
  );
  CEMux inmux_15_17_62460_62528 (
    .I(net_62460),
    .O(net_62528)
  );
  InMux inmux_15_17_62467_62515 (
    .I(net_62467),
    .O(net_62515)
  );
  InMux inmux_15_17_62469_62484 (
    .I(net_62469),
    .O(net_62484)
  );
  InMux inmux_15_17_62470_62488 (
    .I(net_62470),
    .O(net_62488)
  );
  InMux inmux_15_17_62471_62503 (
    .I(net_62471),
    .O(net_62503)
  );
  InMux inmux_15_17_62471_62513 (
    .I(net_62471),
    .O(net_62513)
  );
  InMux inmux_15_17_62472_62490 (
    .I(net_62472),
    .O(net_62490)
  );
  InMux inmux_15_17_62478_62489 (
    .I(net_62478),
    .O(net_62489)
  );
  InMux inmux_15_17_62479_62495 (
    .I(net_62479),
    .O(net_62495)
  );
  ClkMux inmux_15_18_5_62652 (
    .I(net_5),
    .O(net_62652)
  );
  InMux inmux_15_18_62572_62612 (
    .I(net_62572),
    .O(net_62612)
  );
  InMux inmux_15_18_62573_62642 (
    .I(net_62573),
    .O(net_62642)
  );
  InMux inmux_15_18_62574_62605 (
    .I(net_62574),
    .O(net_62605)
  );
  InMux inmux_15_18_62574_62641 (
    .I(net_62574),
    .O(net_62641)
  );
  InMux inmux_15_18_62578_62607 (
    .I(net_62578),
    .O(net_62607)
  );
  InMux inmux_15_18_62579_62644 (
    .I(net_62579),
    .O(net_62644)
  );
  InMux inmux_15_18_62582_62606 (
    .I(net_62582),
    .O(net_62606)
  );
  InMux inmux_15_18_62584_62613 (
    .I(net_62584),
    .O(net_62613)
  );
  InMux inmux_15_18_62588_62614 (
    .I(net_62588),
    .O(net_62614)
  );
  InMux inmux_15_18_62589_62611 (
    .I(net_62589),
    .O(net_62611)
  );
  InMux inmux_15_18_62592_62650 (
    .I(net_62592),
    .O(net_62650)
  );
  InMux inmux_15_18_62593_62632 (
    .I(net_62593),
    .O(net_62632)
  );
  InMux inmux_15_18_62597_62643 (
    .I(net_62597),
    .O(net_62643)
  );
  InMux inmux_15_18_62599_62619 (
    .I(net_62599),
    .O(net_62619)
  );
  InMux inmux_15_18_62600_62608 (
    .I(net_62600),
    .O(net_62608)
  );
  CEMux inmux_15_18_8_62651 (
    .I(net_8),
    .O(net_62651)
  );
  ClkMux inmux_15_19_5_62775 (
    .I(net_5),
    .O(net_62775)
  );
  InMux inmux_15_19_62702_62729 (
    .I(net_62702),
    .O(net_62729)
  );
  InMux inmux_15_19_62703_62748 (
    .I(net_62703),
    .O(net_62748)
  );
  CEMux inmux_15_19_62706_62774 (
    .I(net_62706),
    .O(net_62774)
  );
  InMux inmux_15_19_62715_62761 (
    .I(net_62715),
    .O(net_62761)
  );
  InMux inmux_15_19_62720_62747 (
    .I(net_62720),
    .O(net_62747)
  );
  InMux inmux_15_19_62722_62766 (
    .I(net_62722),
    .O(net_62766)
  );
  InMux inmux_15_19_62723_62746 (
    .I(net_62723),
    .O(net_62746)
  );
  InMux inmux_15_19_62724_62764 (
    .I(net_62724),
    .O(net_62764)
  );
  ClkMux inmux_15_20_5_62898 (
    .I(net_5),
    .O(net_62898)
  );
  InMux inmux_15_20_62818_62851 (
    .I(net_62818),
    .O(net_62851)
  );
  InMux inmux_15_20_62818_62863 (
    .I(net_62818),
    .O(net_62863)
  );
  InMux inmux_15_20_62818_62894 (
    .I(net_62818),
    .O(net_62894)
  );
  InMux inmux_15_20_62821_62888 (
    .I(net_62821),
    .O(net_62888)
  );
  InMux inmux_15_20_62828_62890 (
    .I(net_62828),
    .O(net_62890)
  );
  CEMux inmux_15_20_62829_62897 (
    .I(net_62829),
    .O(net_62897)
  );
  InMux inmux_15_20_62833_62889 (
    .I(net_62833),
    .O(net_62889)
  );
  InMux inmux_15_20_62834_62887 (
    .I(net_62834),
    .O(net_62887)
  );
  SRMux inmux_15_20_62838_62899 (
    .I(net_62838),
    .O(net_62899)
  );
  InMux inmux_15_20_62844_62895 (
    .I(net_62844),
    .O(net_62895)
  );
  InMux inmux_15_20_62849_62865 (
    .I(net_62849),
    .O(net_62865)
  );
  InMux inmux_15_21_62956_63010 (
    .I(net_62956),
    .O(net_63010)
  );
  InMux inmux_15_21_62967_63011 (
    .I(net_62967),
    .O(net_63011)
  );
  ClkMux inmux_15_22_5_63144 (
    .I(net_5),
    .O(net_63144)
  );
  InMux inmux_15_22_63068_63130 (
    .I(net_63068),
    .O(net_63130)
  );
  InMux inmux_15_22_63079_63121 (
    .I(net_63079),
    .O(net_63121)
  );
  CEMux inmux_15_22_63091_63143 (
    .I(net_63091),
    .O(net_63143)
  );
  ClkMux inmux_15_23_5_63267 (
    .I(net_5),
    .O(net_63267)
  );
  InMux inmux_15_23_63191_63251 (
    .I(net_63191),
    .O(net_63251)
  );
  InMux inmux_15_23_63191_63265 (
    .I(net_63191),
    .O(net_63265)
  );
  InMux inmux_15_23_63192_63228 (
    .I(net_63192),
    .O(net_63228)
  );
  InMux inmux_15_23_63192_63252 (
    .I(net_63192),
    .O(net_63252)
  );
  InMux inmux_15_23_63192_63264 (
    .I(net_63192),
    .O(net_63264)
  );
  InMux inmux_15_23_63200_63253 (
    .I(net_63200),
    .O(net_63253)
  );
  InMux inmux_15_23_63200_63263 (
    .I(net_63200),
    .O(net_63263)
  );
  InMux inmux_15_23_63204_63250 (
    .I(net_63204),
    .O(net_63250)
  );
  InMux inmux_15_23_63204_63262 (
    .I(net_63204),
    .O(net_63262)
  );
  CEMux inmux_15_23_63205_63266 (
    .I(net_63205),
    .O(net_63266)
  );
  ClkMux inmux_15_25_5_63513 (
    .I(net_5),
    .O(net_63513)
  );
  InMux inmux_15_25_63439_63499 (
    .I(net_63439),
    .O(net_63499)
  );
  CEMux inmux_15_25_63444_63512 (
    .I(net_63444),
    .O(net_63512)
  );
  InMux inmux_15_27_63683_63743 (
    .I(net_63683),
    .O(net_63743)
  );
  InMux inmux_15_27_63710_63745 (
    .I(net_63710),
    .O(net_63745)
  );
  InMux inmux_15_28_63807_63841 (
    .I(net_63807),
    .O(net_63841)
  );
  InMux inmux_15_28_63819_63838 (
    .I(net_63819),
    .O(net_63838)
  );
  InMux inmux_15_28_63819_63860 (
    .I(net_63819),
    .O(net_63860)
  );
  InMux inmux_15_28_63819_63865 (
    .I(net_63819),
    .O(net_63865)
  );
  InMux inmux_15_28_63819_63879 (
    .I(net_63819),
    .O(net_63879)
  );
  InMux inmux_15_28_63823_63836 (
    .I(net_63823),
    .O(net_63836)
  );
  InMux inmux_15_28_63823_63862 (
    .I(net_63823),
    .O(net_63862)
  );
  InMux inmux_15_28_63823_63877 (
    .I(net_63823),
    .O(net_63877)
  );
  InMux inmux_15_28_63824_63835 (
    .I(net_63824),
    .O(net_63835)
  );
  InMux inmux_15_28_63824_63861 (
    .I(net_63824),
    .O(net_63861)
  );
  InMux inmux_15_28_63824_63868 (
    .I(net_63824),
    .O(net_63868)
  );
  InMux inmux_15_28_63824_63878 (
    .I(net_63824),
    .O(net_63878)
  );
  InMux inmux_15_28_63829_63837 (
    .I(net_63829),
    .O(net_63837)
  );
  InMux inmux_15_28_63829_63842 (
    .I(net_63829),
    .O(net_63842)
  );
  InMux inmux_15_28_63829_63859 (
    .I(net_63829),
    .O(net_63859)
  );
  InMux inmux_15_28_63829_63880 (
    .I(net_63829),
    .O(net_63880)
  );
  InMux inmux_15_28_63830_63867 (
    .I(net_63830),
    .O(net_63867)
  );
  InMux inmux_15_28_63831_63866 (
    .I(net_63831),
    .O(net_63866)
  );
  InMux inmux_15_29_63928_63990 (
    .I(net_63928),
    .O(net_63990)
  );
  InMux inmux_15_29_63930_64002 (
    .I(net_63930),
    .O(net_64002)
  );
  InMux inmux_15_29_63934_63989 (
    .I(net_63934),
    .O(net_63989)
  );
  InMux inmux_15_29_63936_64001 (
    .I(net_63936),
    .O(net_64001)
  );
  InMux inmux_15_29_63938_63991 (
    .I(net_63938),
    .O(net_63991)
  );
  InMux inmux_15_29_63939_63988 (
    .I(net_63939),
    .O(net_63988)
  );
  InMux inmux_15_29_63954_64003 (
    .I(net_63954),
    .O(net_64003)
  );
  ClkMux inmux_15_2_5_60684 (
    .I(net_5),
    .O(net_60684)
  );
  InMux inmux_15_2_60604_60639 (
    .I(net_60604),
    .O(net_60639)
  );
  InMux inmux_15_2_60604_60644 (
    .I(net_60604),
    .O(net_60644)
  );
  InMux inmux_15_2_60604_60651 (
    .I(net_60604),
    .O(net_60651)
  );
  InMux inmux_15_2_60604_60656 (
    .I(net_60604),
    .O(net_60656)
  );
  CEMux inmux_15_2_60606_60683 (
    .I(net_60606),
    .O(net_60683)
  );
  InMux inmux_15_2_60610_60637 (
    .I(net_60610),
    .O(net_60637)
  );
  InMux inmux_15_2_60610_60649 (
    .I(net_60610),
    .O(net_60649)
  );
  InMux inmux_15_2_60611_60638 (
    .I(net_60611),
    .O(net_60638)
  );
  InMux inmux_15_2_60611_60645 (
    .I(net_60611),
    .O(net_60645)
  );
  InMux inmux_15_2_60611_60650 (
    .I(net_60611),
    .O(net_60650)
  );
  InMux inmux_15_2_60611_60657 (
    .I(net_60611),
    .O(net_60657)
  );
  InMux inmux_15_2_60614_60643 (
    .I(net_60614),
    .O(net_60643)
  );
  InMux inmux_15_2_60614_60655 (
    .I(net_60614),
    .O(net_60655)
  );
  InMux inmux_15_2_60614_60676 (
    .I(net_60614),
    .O(net_60676)
  );
  InMux inmux_15_2_60615_60646 (
    .I(net_60615),
    .O(net_60646)
  );
  InMux inmux_15_2_60615_60658 (
    .I(net_60615),
    .O(net_60658)
  );
  InMux inmux_15_2_60615_60673 (
    .I(net_60615),
    .O(net_60673)
  );
  InMux inmux_15_2_60628_60652 (
    .I(net_60628),
    .O(net_60652)
  );
  ClkMux inmux_15_3_5_60807 (
    .I(net_5),
    .O(net_60807)
  );
  CEMux inmux_15_3_60729_60806 (
    .I(net_60729),
    .O(net_60806)
  );
  InMux inmux_15_3_60732_60787 (
    .I(net_60732),
    .O(net_60787)
  );
  InMux inmux_15_3_60735_60792 (
    .I(net_60735),
    .O(net_60792)
  );
  InMux inmux_15_3_60735_60797 (
    .I(net_60735),
    .O(net_60797)
  );
  InMux inmux_15_3_60735_60804 (
    .I(net_60735),
    .O(net_60804)
  );
  InMux inmux_15_3_60736_60793 (
    .I(net_60736),
    .O(net_60793)
  );
  InMux inmux_15_3_60738_60769 (
    .I(net_60738),
    .O(net_60769)
  );
  InMux inmux_15_3_60738_60786 (
    .I(net_60738),
    .O(net_60786)
  );
  InMux inmux_15_3_60738_60796 (
    .I(net_60738),
    .O(net_60796)
  );
  InMux inmux_15_3_60738_60805 (
    .I(net_60738),
    .O(net_60805)
  );
  InMux inmux_15_3_60739_60773 (
    .I(net_60739),
    .O(net_60773)
  );
  InMux inmux_15_3_60739_60778 (
    .I(net_60739),
    .O(net_60778)
  );
  InMux inmux_15_3_60740_60781 (
    .I(net_60740),
    .O(net_60781)
  );
  InMux inmux_15_3_60740_60784 (
    .I(net_60740),
    .O(net_60784)
  );
  InMux inmux_15_3_60747_60772 (
    .I(net_60747),
    .O(net_60772)
  );
  InMux inmux_15_3_60749_60779 (
    .I(net_60749),
    .O(net_60779)
  );
  InMux inmux_15_3_60753_60768 (
    .I(net_60753),
    .O(net_60768)
  );
  InMux inmux_15_3_60753_60785 (
    .I(net_60753),
    .O(net_60785)
  );
  InMux inmux_15_3_60753_60799 (
    .I(net_60753),
    .O(net_60799)
  );
  InMux inmux_15_3_60753_60802 (
    .I(net_60753),
    .O(net_60802)
  );
  InMux inmux_15_3_60754_60767 (
    .I(net_60754),
    .O(net_60767)
  );
  InMux inmux_15_3_60758_60791 (
    .I(net_60758),
    .O(net_60791)
  );
  InMux inmux_15_3_60758_60798 (
    .I(net_60758),
    .O(net_60798)
  );
  InMux inmux_15_3_60758_60803 (
    .I(net_60758),
    .O(net_60803)
  );
  ClkMux inmux_15_6_5_61176 (
    .I(net_5),
    .O(net_61176)
  );
  InMux inmux_15_6_61119_61144 (
    .I(net_61119),
    .O(net_61144)
  );
  CEMux inmux_15_6_61123_61175 (
    .I(net_61123),
    .O(net_61175)
  );
  ClkMux inmux_15_8_5_61422 (
    .I(net_5),
    .O(net_61422)
  );
  InMux inmux_15_8_61350_61376 (
    .I(net_61350),
    .O(net_61376)
  );
  CEMux inmux_15_8_61353_61421 (
    .I(net_61353),
    .O(net_61421)
  );
  ClkMux inmux_15_9_5_61545 (
    .I(net_5),
    .O(net_61545)
  );
  InMux inmux_15_9_61473_61540 (
    .I(net_61473),
    .O(net_61540)
  );
  CEMux inmux_15_9_61476_61544 (
    .I(net_61476),
    .O(net_61544)
  );
  InMux inmux_15_9_61483_61498 (
    .I(net_61483),
    .O(net_61498)
  );
  SRMux inmux_15_9_61485_61546 (
    .I(net_61485),
    .O(net_61546)
  );
  InMux inmux_15_9_61486_61501 (
    .I(net_61486),
    .O(net_61501)
  );
  InMux inmux_15_9_61486_61530 (
    .I(net_61486),
    .O(net_61530)
  );
  InMux inmux_15_9_61486_61542 (
    .I(net_61486),
    .O(net_61542)
  );
  InMux inmux_16_10_65428_65485 (
    .I(net_65428),
    .O(net_65485)
  );
  ClkMux inmux_16_11_5_65622 (
    .I(net_5),
    .O(net_65622)
  );
  InMux inmux_16_11_65547_65600 (
    .I(net_65547),
    .O(net_65600)
  );
  InMux inmux_16_11_65548_65608 (
    .I(net_65548),
    .O(net_65608)
  );
  InMux inmux_16_11_65552_65576 (
    .I(net_65552),
    .O(net_65576)
  );
  InMux inmux_16_11_65566_65583 (
    .I(net_65566),
    .O(net_65583)
  );
  CEMux inmux_16_11_8_65621 (
    .I(net_8),
    .O(net_65621)
  );
  ClkMux inmux_16_12_5_65745 (
    .I(net_5),
    .O(net_65745)
  );
  InMux inmux_16_12_65667_65707 (
    .I(net_65667),
    .O(net_65707)
  );
  InMux inmux_16_12_65674_65698 (
    .I(net_65674),
    .O(net_65698)
  );
  InMux inmux_16_12_65674_65705 (
    .I(net_65674),
    .O(net_65705)
  );
  InMux inmux_16_12_65674_65729 (
    .I(net_65674),
    .O(net_65729)
  );
  InMux inmux_16_12_65674_65736 (
    .I(net_65674),
    .O(net_65736)
  );
  InMux inmux_16_12_65675_65730 (
    .I(net_65675),
    .O(net_65730)
  );
  InMux inmux_16_12_65677_65701 (
    .I(net_65677),
    .O(net_65701)
  );
  InMux inmux_16_12_65678_65734 (
    .I(net_65678),
    .O(net_65734)
  );
  InMux inmux_16_12_65679_65737 (
    .I(net_65679),
    .O(net_65737)
  );
  InMux inmux_16_12_65680_65712 (
    .I(net_65680),
    .O(net_65712)
  );
  InMux inmux_16_12_65683_65731 (
    .I(net_65683),
    .O(net_65731)
  );
  InMux inmux_16_12_65684_65699 (
    .I(net_65684),
    .O(net_65699)
  );
  InMux inmux_16_12_65686_65706 (
    .I(net_65686),
    .O(net_65706)
  );
  InMux inmux_16_12_65687_65700 (
    .I(net_65687),
    .O(net_65700)
  );
  InMux inmux_16_12_65688_65735 (
    .I(net_65688),
    .O(net_65735)
  );
  InMux inmux_16_12_65689_65728 (
    .I(net_65689),
    .O(net_65728)
  );
  InMux inmux_16_12_65693_65704 (
    .I(net_65693),
    .O(net_65704)
  );
  InMux inmux_16_12_65695_65723 (
    .I(net_65695),
    .O(net_65723)
  );
  CEMux inmux_16_12_8_65744 (
    .I(net_8),
    .O(net_65744)
  );
  ClkMux inmux_16_13_5_65868 (
    .I(net_5),
    .O(net_65868)
  );
  InMux inmux_16_13_65790_65821 (
    .I(net_65790),
    .O(net_65821)
  );
  InMux inmux_16_13_65791_65836 (
    .I(net_65791),
    .O(net_65836)
  );
  InMux inmux_16_13_65792_65833 (
    .I(net_65792),
    .O(net_65833)
  );
  InMux inmux_16_13_65801_65835 (
    .I(net_65801),
    .O(net_65835)
  );
  InMux inmux_16_13_65806_65842 (
    .I(net_65806),
    .O(net_65842)
  );
  InMux inmux_16_13_65807_65834 (
    .I(net_65807),
    .O(net_65834)
  );
  InMux inmux_16_13_65812_65846 (
    .I(net_65812),
    .O(net_65846)
  );
  InMux inmux_16_13_65814_65848 (
    .I(net_65814),
    .O(net_65848)
  );
  ClkMux inmux_16_14_5_65991 (
    .I(net_5),
    .O(net_65991)
  );
  InMux inmux_16_14_65917_65987 (
    .I(net_65917),
    .O(net_65987)
  );
  InMux inmux_16_14_65918_65976 (
    .I(net_65918),
    .O(net_65976)
  );
  InMux inmux_16_14_65935_65974 (
    .I(net_65935),
    .O(net_65974)
  );
  InMux inmux_16_14_65937_65952 (
    .I(net_65937),
    .O(net_65952)
  );
  InMux inmux_16_14_65942_65953 (
    .I(net_65942),
    .O(net_65953)
  );
  CEMux inmux_16_14_6_65990 (
    .I(net_6),
    .O(net_65990)
  );
  ClkMux inmux_16_15_5_66114 (
    .I(net_5),
    .O(net_66114)
  );
  InMux inmux_16_15_66034_66110 (
    .I(net_66034),
    .O(net_66110)
  );
  InMux inmux_16_15_66035_66097 (
    .I(net_66035),
    .O(net_66097)
  );
  InMux inmux_16_15_66036_66069 (
    .I(net_66036),
    .O(net_66069)
  );
  InMux inmux_16_15_66040_66103 (
    .I(net_66040),
    .O(net_66103)
  );
  InMux inmux_16_15_66041_66106 (
    .I(net_66041),
    .O(net_66106)
  );
  InMux inmux_16_15_66042_66068 (
    .I(net_66042),
    .O(net_66068)
  );
  InMux inmux_16_15_66042_66085 (
    .I(net_66042),
    .O(net_66085)
  );
  InMux inmux_16_15_66042_66094 (
    .I(net_66042),
    .O(net_66094)
  );
  InMux inmux_16_15_66042_66099 (
    .I(net_66042),
    .O(net_66099)
  );
  InMux inmux_16_15_66049_66098 (
    .I(net_66049),
    .O(net_66098)
  );
  InMux inmux_16_15_66050_66079 (
    .I(net_66050),
    .O(net_66079)
  );
  InMux inmux_16_15_66054_66091 (
    .I(net_66054),
    .O(net_66091)
  );
  InMux inmux_16_15_66055_66080 (
    .I(net_66055),
    .O(net_66080)
  );
  InMux inmux_16_15_66056_66100 (
    .I(net_66056),
    .O(net_66100)
  );
  InMux inmux_16_15_66057_66082 (
    .I(net_66057),
    .O(net_66082)
  );
  InMux inmux_16_15_66057_66104 (
    .I(net_66057),
    .O(net_66104)
  );
  InMux inmux_16_15_66061_66105 (
    .I(net_66061),
    .O(net_66105)
  );
  InMux inmux_16_15_66062_66087 (
    .I(net_66062),
    .O(net_66087)
  );
  InMux inmux_16_15_66065_66081 (
    .I(net_66065),
    .O(net_66081)
  );
  CEMux inmux_16_15_8_66113 (
    .I(net_8),
    .O(net_66113)
  );
  ClkMux inmux_16_16_5_66237 (
    .I(net_5),
    .O(net_66237)
  );
  InMux inmux_16_16_66158_66198 (
    .I(net_66158),
    .O(net_66198)
  );
  InMux inmux_16_16_66178_66203 (
    .I(net_66178),
    .O(net_66203)
  );
  InMux inmux_16_16_66181_66196 (
    .I(net_66181),
    .O(net_66196)
  );
  CEMux inmux_16_16_66184_66236 (
    .I(net_66184),
    .O(net_66236)
  );
  CEMux inmux_16_17_10_66359 (
    .I(net_10),
    .O(net_66359)
  );
  ClkMux inmux_16_17_5_66360 (
    .I(net_5),
    .O(net_66360)
  );
  InMux inmux_16_17_66281_66321 (
    .I(net_66281),
    .O(net_66321)
  );
  ClkMux inmux_16_18_5_66483 (
    .I(net_5),
    .O(net_66483)
  );
  InMux inmux_16_18_66405_66448 (
    .I(net_66405),
    .O(net_66448)
  );
  InMux inmux_16_18_66408_66451 (
    .I(net_66408),
    .O(net_66451)
  );
  CEMux inmux_16_18_66414_66482 (
    .I(net_66414),
    .O(net_66482)
  );
  InMux inmux_16_18_66415_66449 (
    .I(net_66415),
    .O(net_66449)
  );
  InMux inmux_16_18_66416_66450 (
    .I(net_66416),
    .O(net_66450)
  );
  InMux inmux_16_18_66422_66463 (
    .I(net_66422),
    .O(net_66463)
  );
  InMux inmux_16_18_66430_66460 (
    .I(net_66430),
    .O(net_66460)
  );
  InMux inmux_16_18_66433_66456 (
    .I(net_66433),
    .O(net_66456)
  );
  ClkMux inmux_16_19_5_66606 (
    .I(net_5),
    .O(net_66606)
  );
  InMux inmux_16_19_66527_66577 (
    .I(net_66527),
    .O(net_66577)
  );
  InMux inmux_16_19_66528_66568 (
    .I(net_66528),
    .O(net_66568)
  );
  InMux inmux_16_19_66531_66596 (
    .I(net_66531),
    .O(net_66596)
  );
  InMux inmux_16_19_66533_66591 (
    .I(net_66533),
    .O(net_66591)
  );
  InMux inmux_16_19_66537_66592 (
    .I(net_66537),
    .O(net_66592)
  );
  InMux inmux_16_19_66538_66565 (
    .I(net_66538),
    .O(net_66565)
  );
  InMux inmux_16_19_66538_66589 (
    .I(net_66538),
    .O(net_66589)
  );
  InMux inmux_16_19_66543_66601 (
    .I(net_66543),
    .O(net_66601)
  );
  InMux inmux_16_19_66546_66566 (
    .I(net_66546),
    .O(net_66566)
  );
  InMux inmux_16_19_66546_66590 (
    .I(net_66546),
    .O(net_66590)
  );
  InMux inmux_16_19_66553_66585 (
    .I(net_66553),
    .O(net_66585)
  );
  InMux inmux_16_19_66554_66567 (
    .I(net_66554),
    .O(net_66567)
  );
  InMux inmux_16_19_66557_66597 (
    .I(net_66557),
    .O(net_66597)
  );
  CEMux inmux_16_19_6_66605 (
    .I(net_6),
    .O(net_66605)
  );
  ClkMux inmux_16_20_5_66729 (
    .I(net_5),
    .O(net_66729)
  );
  InMux inmux_16_20_66650_66700 (
    .I(net_66650),
    .O(net_66700)
  );
  InMux inmux_16_20_66650_66714 (
    .I(net_66650),
    .O(net_66714)
  );
  InMux inmux_16_20_66652_66690 (
    .I(net_66652),
    .O(net_66690)
  );
  InMux inmux_16_20_66653_66715 (
    .I(net_66653),
    .O(net_66715)
  );
  InMux inmux_16_20_66656_66712 (
    .I(net_66656),
    .O(net_66712)
  );
  InMux inmux_16_20_66658_66713 (
    .I(net_66658),
    .O(net_66713)
  );
  CEMux inmux_16_20_66660_66728 (
    .I(net_66660),
    .O(net_66728)
  );
  InMux inmux_16_20_66661_66724 (
    .I(net_66661),
    .O(net_66724)
  );
  InMux inmux_16_20_66664_66701 (
    .I(net_66664),
    .O(net_66701)
  );
  InMux inmux_16_20_66667_66708 (
    .I(net_66667),
    .O(net_66708)
  );
  InMux inmux_16_20_66674_66703 (
    .I(net_66674),
    .O(net_66703)
  );
  InMux inmux_16_20_66675_66702 (
    .I(net_66675),
    .O(net_66702)
  );
  InMux inmux_16_20_66676_66696 (
    .I(net_66676),
    .O(net_66696)
  );
  ClkMux inmux_16_21_5_66852 (
    .I(net_5),
    .O(net_66852)
  );
  InMux inmux_16_21_66797_66850 (
    .I(net_66797),
    .O(net_66850)
  );
  CEMux inmux_16_21_6_66851 (
    .I(net_6),
    .O(net_66851)
  );
  ClkMux inmux_16_28_5_67713 (
    .I(net_5),
    .O(net_67713)
  );
  InMux inmux_16_28_67633_67704 (
    .I(net_67633),
    .O(net_67704)
  );
  CEMux inmux_16_28_67635_67712 (
    .I(net_67635),
    .O(net_67712)
  );
  InMux inmux_16_28_67637_67675 (
    .I(net_67637),
    .O(net_67675)
  );
  InMux inmux_16_28_67637_67678 (
    .I(net_67637),
    .O(net_67678)
  );
  InMux inmux_16_28_67642_67685 (
    .I(net_67642),
    .O(net_67685)
  );
  InMux inmux_16_28_67642_67697 (
    .I(net_67642),
    .O(net_67697)
  );
  InMux inmux_16_28_67642_67711 (
    .I(net_67642),
    .O(net_67711)
  );
  InMux inmux_16_28_67643_67674 (
    .I(net_67643),
    .O(net_67674)
  );
  InMux inmux_16_28_67645_67681 (
    .I(net_67645),
    .O(net_67681)
  );
  InMux inmux_16_28_67647_67686 (
    .I(net_67647),
    .O(net_67686)
  );
  InMux inmux_16_28_67647_67698 (
    .I(net_67647),
    .O(net_67698)
  );
  InMux inmux_16_28_67647_67705 (
    .I(net_67647),
    .O(net_67705)
  );
  InMux inmux_16_28_67647_67710 (
    .I(net_67647),
    .O(net_67710)
  );
  InMux inmux_16_28_67649_67673 (
    .I(net_67649),
    .O(net_67673)
  );
  InMux inmux_16_28_67649_67702 (
    .I(net_67649),
    .O(net_67702)
  );
  InMux inmux_16_28_67650_67672 (
    .I(net_67650),
    .O(net_67672)
  );
  InMux inmux_16_28_67650_67703 (
    .I(net_67650),
    .O(net_67703)
  );
  InMux inmux_16_28_67654_67679 (
    .I(net_67654),
    .O(net_67679)
  );
  InMux inmux_16_28_67654_67684 (
    .I(net_67654),
    .O(net_67684)
  );
  InMux inmux_16_28_67654_67696 (
    .I(net_67654),
    .O(net_67696)
  );
  InMux inmux_16_28_67654_67708 (
    .I(net_67654),
    .O(net_67708)
  );
  InMux inmux_16_28_67656_67693 (
    .I(net_67656),
    .O(net_67693)
  );
  InMux inmux_16_28_67657_67691 (
    .I(net_67657),
    .O(net_67691)
  );
  InMux inmux_16_28_67660_67680 (
    .I(net_67660),
    .O(net_67680)
  );
  InMux inmux_16_28_67660_67687 (
    .I(net_67660),
    .O(net_67687)
  );
  InMux inmux_16_28_67660_67699 (
    .I(net_67660),
    .O(net_67699)
  );
  InMux inmux_16_28_67660_67709 (
    .I(net_67660),
    .O(net_67709)
  );
  ClkMux inmux_16_29_5_67836 (
    .I(net_5),
    .O(net_67836)
  );
  InMux inmux_16_29_67757_67790 (
    .I(net_67757),
    .O(net_67790)
  );
  CEMux inmux_16_29_67758_67835 (
    .I(net_67758),
    .O(net_67835)
  );
  InMux inmux_16_29_67759_67802 (
    .I(net_67759),
    .O(net_67802)
  );
  InMux inmux_16_29_67759_67816 (
    .I(net_67759),
    .O(net_67816)
  );
  InMux inmux_16_29_67761_67792 (
    .I(net_67761),
    .O(net_67792)
  );
  InMux inmux_16_29_67765_67815 (
    .I(net_67765),
    .O(net_67815)
  );
  InMux inmux_16_29_67767_67791 (
    .I(net_67767),
    .O(net_67791)
  );
  InMux inmux_16_29_67770_67814 (
    .I(net_67770),
    .O(net_67814)
  );
  InMux inmux_16_29_67772_67825 (
    .I(net_67772),
    .O(net_67825)
  );
  InMux inmux_16_29_67774_67813 (
    .I(net_67774),
    .O(net_67813)
  );
  InMux inmux_16_29_67774_67827 (
    .I(net_67774),
    .O(net_67827)
  );
  InMux inmux_16_29_67778_67789 (
    .I(net_67778),
    .O(net_67789)
  );
  ClkMux inmux_16_2_5_64515 (
    .I(net_5),
    .O(net_64515)
  );
  InMux inmux_16_2_64436_64488 (
    .I(net_64436),
    .O(net_64488)
  );
  InMux inmux_16_2_64443_64483 (
    .I(net_64443),
    .O(net_64483)
  );
  InMux inmux_16_2_64443_64500 (
    .I(net_64443),
    .O(net_64500)
  );
  InMux inmux_16_2_64444_64499 (
    .I(net_64444),
    .O(net_64499)
  );
  InMux inmux_16_2_64449_64481 (
    .I(net_64449),
    .O(net_64481)
  );
  InMux inmux_16_2_64455_64475 (
    .I(net_64455),
    .O(net_64475)
  );
  InMux inmux_16_2_64455_64501 (
    .I(net_64455),
    .O(net_64501)
  );
  InMux inmux_16_2_64458_64498 (
    .I(net_64458),
    .O(net_64498)
  );
  InMux inmux_16_2_64461_64486 (
    .I(net_64461),
    .O(net_64486)
  );
  CEMux inmux_16_2_64462_64514 (
    .I(net_64462),
    .O(net_64514)
  );
  InMux inmux_16_2_64466_64480 (
    .I(net_64466),
    .O(net_64480)
  );
  InMux inmux_16_5_64814_64838 (
    .I(net_64814),
    .O(net_64838)
  );
  InMux inmux_16_5_64818_64845 (
    .I(net_64818),
    .O(net_64845)
  );
  InMux inmux_16_5_64820_64856 (
    .I(net_64820),
    .O(net_64856)
  );
  InMux inmux_16_5_64827_64874 (
    .I(net_64827),
    .O(net_64874)
  );
  InMux inmux_16_5_64829_64880 (
    .I(net_64829),
    .O(net_64880)
  );
  InMux inmux_16_5_64830_64850 (
    .I(net_64830),
    .O(net_64850)
  );
  InMux inmux_16_5_64831_64868 (
    .I(net_64831),
    .O(net_64868)
  );
  InMux inmux_16_5_64834_64862 (
    .I(net_64834),
    .O(net_64862)
  );
  InMux inmux_16_5_64842_64852 (
    .I(net_64842),
    .O(net_64852)
  );
  InMux inmux_16_5_64848_64858 (
    .I(net_64848),
    .O(net_64858)
  );
  InMux inmux_16_5_64854_64864 (
    .I(net_64854),
    .O(net_64864)
  );
  InMux inmux_16_5_64860_64870 (
    .I(net_64860),
    .O(net_64870)
  );
  InMux inmux_16_5_64866_64876 (
    .I(net_64866),
    .O(net_64876)
  );
  InMux inmux_16_5_64872_64882 (
    .I(net_64872),
    .O(net_64882)
  );
  InMux inmux_16_6_64922_64963 (
    .I(net_64922),
    .O(net_64963)
  );
  InMux inmux_16_6_64943_64962 (
    .I(net_64943),
    .O(net_64962)
  );
  ClkMux inmux_16_9_5_65376 (
    .I(net_5),
    .O(net_65376)
  );
  InMux inmux_16_9_65298_65372 (
    .I(net_65298),
    .O(net_65372)
  );
  InMux inmux_16_9_65302_65355 (
    .I(net_65302),
    .O(net_65355)
  );
  InMux inmux_16_9_65304_65371 (
    .I(net_65304),
    .O(net_65371)
  );
  CEMux inmux_16_9_65307_65375 (
    .I(net_65307),
    .O(net_65375)
  );
  InMux inmux_16_9_65308_65342 (
    .I(net_65308),
    .O(net_65342)
  );
  InMux inmux_16_9_65308_65361 (
    .I(net_65308),
    .O(net_65361)
  );
  InMux inmux_16_9_65315_65344 (
    .I(net_65315),
    .O(net_65344)
  );
  InMux inmux_16_9_65315_65359 (
    .I(net_65315),
    .O(net_65359)
  );
  InMux inmux_16_9_65318_65343 (
    .I(net_65318),
    .O(net_65343)
  );
  InMux inmux_16_9_65318_65350 (
    .I(net_65318),
    .O(net_65350)
  );
  InMux inmux_16_9_65318_65362 (
    .I(net_65318),
    .O(net_65362)
  );
  InMux inmux_16_9_65321_65341 (
    .I(net_65321),
    .O(net_65341)
  );
  InMux inmux_16_9_65321_65360 (
    .I(net_65321),
    .O(net_65360)
  );
  InMux inmux_16_9_65321_65367 (
    .I(net_65321),
    .O(net_65367)
  );
  ClkMux inmux_17_0_5_68043 (
    .I(net_5),
    .O(net_68043)
  );
  ClkMux inmux_17_0_5_68044 (
    .I(net_5),
    .O(net_68044)
  );
  IoInMux inmux_17_0_68056_68036 (
    .I(net_68056),
    .O(net_68036)
  );
  CEMux inmux_17_0_68058_68042 (
    .I(net_68058),
    .O(net_68042)
  );
  ClkMux inmux_17_12_5_69576 (
    .I(net_5),
    .O(net_69576)
  );
  InMux inmux_17_12_69503_69535 (
    .I(net_69503),
    .O(net_69535)
  );
  SRMux inmux_17_12_69525_69577 (
    .I(net_69525),
    .O(net_69577)
  );
  CEMux inmux_17_13_10_69698 (
    .I(net_10),
    .O(net_69698)
  );
  SRMux inmux_17_13_11_69700 (
    .I(net_11),
    .O(net_69700)
  );
  ClkMux inmux_17_13_5_69699 (
    .I(net_5),
    .O(net_69699)
  );
  InMux inmux_17_13_69619_69690 (
    .I(net_69619),
    .O(net_69690)
  );
  InMux inmux_17_13_69623_69671 (
    .I(net_69623),
    .O(net_69671)
  );
  InMux inmux_17_13_69627_69689 (
    .I(net_69627),
    .O(net_69689)
  );
  InMux inmux_17_13_69629_69670 (
    .I(net_69629),
    .O(net_69670)
  );
  InMux inmux_17_13_69629_69691 (
    .I(net_69629),
    .O(net_69691)
  );
  InMux inmux_17_13_69630_69673 (
    .I(net_69630),
    .O(net_69673)
  );
  ClkMux inmux_17_14_5_69822 (
    .I(net_5),
    .O(net_69822)
  );
  InMux inmux_17_14_69742_69806 (
    .I(net_69742),
    .O(net_69806)
  );
  InMux inmux_17_14_69747_69788 (
    .I(net_69747),
    .O(net_69788)
  );
  InMux inmux_17_14_69749_69807 (
    .I(net_69749),
    .O(net_69807)
  );
  InMux inmux_17_14_69750_69802 (
    .I(net_69750),
    .O(net_69802)
  );
  InMux inmux_17_14_69753_69808 (
    .I(net_69753),
    .O(net_69808)
  );
  InMux inmux_17_14_69754_69805 (
    .I(net_69754),
    .O(net_69805)
  );
  InMux inmux_17_14_69756_69778 (
    .I(net_69756),
    .O(net_69778)
  );
  InMux inmux_17_14_69760_69796 (
    .I(net_69760),
    .O(net_69796)
  );
  InMux inmux_17_14_69763_69817 (
    .I(net_69763),
    .O(net_69817)
  );
  CEMux inmux_17_15_10_69944 (
    .I(net_10),
    .O(net_69944)
  );
  SRMux inmux_17_15_11_69946 (
    .I(net_11),
    .O(net_69946)
  );
  ClkMux inmux_17_15_5_69945 (
    .I(net_5),
    .O(net_69945)
  );
  InMux inmux_17_15_69865_69924 (
    .I(net_69865),
    .O(net_69924)
  );
  InMux inmux_17_15_69867_69900 (
    .I(net_69867),
    .O(net_69900)
  );
  InMux inmux_17_15_69873_69923 (
    .I(net_69873),
    .O(net_69923)
  );
  InMux inmux_17_15_69875_69925 (
    .I(net_69875),
    .O(net_69925)
  );
  InMux inmux_17_15_69877_69918 (
    .I(net_69877),
    .O(net_69918)
  );
  InMux inmux_17_15_69878_69919 (
    .I(net_69878),
    .O(net_69919)
  );
  InMux inmux_17_15_69879_69916 (
    .I(net_69879),
    .O(net_69916)
  );
  InMux inmux_17_15_69880_69898 (
    .I(net_69880),
    .O(net_69898)
  );
  ClkMux inmux_17_16_5_70068 (
    .I(net_5),
    .O(net_70068)
  );
  InMux inmux_17_16_70003_70030 (
    .I(net_70003),
    .O(net_70030)
  );
  InMux inmux_17_16_70014_70065 (
    .I(net_70014),
    .O(net_70065)
  );
  SRMux inmux_17_16_70017_70069 (
    .I(net_70017),
    .O(net_70069)
  );
  CEMux inmux_17_17_10_70190 (
    .I(net_10),
    .O(net_70190)
  );
  SRMux inmux_17_17_11_70192 (
    .I(net_11),
    .O(net_70192)
  );
  ClkMux inmux_17_17_5_70191 (
    .I(net_5),
    .O(net_70191)
  );
  InMux inmux_17_17_70112_70145 (
    .I(net_70112),
    .O(net_70145)
  );
  InMux inmux_17_17_70113_70156 (
    .I(net_70113),
    .O(net_70156)
  );
  InMux inmux_17_17_70120_70187 (
    .I(net_70120),
    .O(net_70187)
  );
  InMux inmux_17_17_70121_70150 (
    .I(net_70121),
    .O(net_70150)
  );
  InMux inmux_17_17_70121_70176 (
    .I(net_70121),
    .O(net_70176)
  );
  InMux inmux_17_17_70123_70188 (
    .I(net_70123),
    .O(net_70188)
  );
  InMux inmux_17_17_70124_70175 (
    .I(net_70124),
    .O(net_70175)
  );
  InMux inmux_17_17_70128_70147 (
    .I(net_70128),
    .O(net_70147)
  );
  InMux inmux_17_17_70128_70157 (
    .I(net_70128),
    .O(net_70157)
  );
  InMux inmux_17_17_70136_70151 (
    .I(net_70136),
    .O(net_70151)
  );
  InMux inmux_17_17_70137_70186 (
    .I(net_70137),
    .O(net_70186)
  );
  InMux inmux_17_17_70138_70158 (
    .I(net_70138),
    .O(net_70158)
  );
  InMux inmux_17_17_70140_70146 (
    .I(net_70140),
    .O(net_70146)
  );
  ClkMux inmux_17_18_5_70314 (
    .I(net_5),
    .O(net_70314)
  );
  InMux inmux_17_18_70236_70288 (
    .I(net_70236),
    .O(net_70288)
  );
  InMux inmux_17_18_70239_70282 (
    .I(net_70239),
    .O(net_70282)
  );
  InMux inmux_17_18_70243_70305 (
    .I(net_70243),
    .O(net_70305)
  );
  InMux inmux_17_18_70245_70269 (
    .I(net_70245),
    .O(net_70269)
  );
  InMux inmux_17_18_70247_70293 (
    .I(net_70247),
    .O(net_70293)
  );
  InMux inmux_17_18_70248_70309 (
    .I(net_70248),
    .O(net_70309)
  );
  InMux inmux_17_18_70254_70274 (
    .I(net_70254),
    .O(net_70274)
  );
  ClkMux inmux_17_19_5_70437 (
    .I(net_5),
    .O(net_70437)
  );
  InMux inmux_17_19_70358_70427 (
    .I(net_70358),
    .O(net_70427)
  );
  InMux inmux_17_19_70362_70417 (
    .I(net_70362),
    .O(net_70417)
  );
  InMux inmux_17_19_70363_70414 (
    .I(net_70363),
    .O(net_70414)
  );
  InMux inmux_17_19_70365_70429 (
    .I(net_70365),
    .O(net_70429)
  );
  InMux inmux_17_19_70371_70398 (
    .I(net_70371),
    .O(net_70398)
  );
  InMux inmux_17_19_70374_70434 (
    .I(net_70374),
    .O(net_70434)
  );
  CEMux inmux_17_19_70375_70436 (
    .I(net_70375),
    .O(net_70436)
  );
  InMux inmux_17_19_70376_70415 (
    .I(net_70376),
    .O(net_70415)
  );
  InMux inmux_17_19_70379_70416 (
    .I(net_70379),
    .O(net_70416)
  );
  InMux inmux_17_19_70379_70433 (
    .I(net_70379),
    .O(net_70433)
  );
  InMux inmux_17_19_70382_70428 (
    .I(net_70382),
    .O(net_70428)
  );
  InMux inmux_17_19_70385_70420 (
    .I(net_70385),
    .O(net_70420)
  );
  InMux inmux_17_19_70388_70426 (
    .I(net_70388),
    .O(net_70426)
  );
  ClkMux inmux_17_20_5_70560 (
    .I(net_5),
    .O(net_70560)
  );
  InMux inmux_17_20_70489_70549 (
    .I(net_70489),
    .O(net_70549)
  );
  InMux inmux_17_20_70493_70520 (
    .I(net_70493),
    .O(net_70520)
  );
  InMux inmux_17_20_70494_70550 (
    .I(net_70494),
    .O(net_70550)
  );
  InMux inmux_17_20_70497_70528 (
    .I(net_70497),
    .O(net_70528)
  );
  InMux inmux_17_20_70501_70519 (
    .I(net_70501),
    .O(net_70519)
  );
  InMux inmux_17_20_70502_70522 (
    .I(net_70502),
    .O(net_70522)
  );
  InMux inmux_17_20_70503_70543 (
    .I(net_70503),
    .O(net_70543)
  );
  InMux inmux_17_20_70507_70515 (
    .I(net_70507),
    .O(net_70515)
  );
  InMux inmux_17_20_70508_70521 (
    .I(net_70508),
    .O(net_70521)
  );
  CEMux inmux_17_20_8_70559 (
    .I(net_8),
    .O(net_70559)
  );
  ClkMux inmux_17_21_5_70683 (
    .I(net_5),
    .O(net_70683)
  );
  CEMux inmux_17_21_70605_70682 (
    .I(net_70605),
    .O(net_70682)
  );
  InMux inmux_17_21_70606_70668 (
    .I(net_70606),
    .O(net_70668)
  );
  InMux inmux_17_21_70620_70675 (
    .I(net_70620),
    .O(net_70675)
  );
  InMux inmux_17_29_71604_71650 (
    .I(net_71604),
    .O(net_71650)
  );
  InMux inmux_17_29_71604_71659 (
    .I(net_71604),
    .O(net_71659)
  );
  InMux inmux_17_29_71604_71664 (
    .I(net_71604),
    .O(net_71664)
  );
  InMux inmux_17_29_71608_71652 (
    .I(net_71608),
    .O(net_71652)
  );
  InMux inmux_17_29_71608_71657 (
    .I(net_71608),
    .O(net_71657)
  );
  InMux inmux_17_29_71608_71662 (
    .I(net_71608),
    .O(net_71662)
  );
  InMux inmux_17_29_71609_71651 (
    .I(net_71609),
    .O(net_71651)
  );
  InMux inmux_17_29_71609_71656 (
    .I(net_71609),
    .O(net_71656)
  );
  InMux inmux_17_29_71609_71663 (
    .I(net_71609),
    .O(net_71663)
  );
  InMux inmux_17_29_71614_71653 (
    .I(net_71614),
    .O(net_71653)
  );
  InMux inmux_17_29_71614_71658 (
    .I(net_71614),
    .O(net_71658)
  );
  InMux inmux_17_29_71614_71665 (
    .I(net_71614),
    .O(net_71665)
  );
  ClkMux inmux_17_31_5_71844 (
    .I(net_5),
    .O(net_71844)
  );
  ClkMux inmux_17_31_5_71845 (
    .I(net_5),
    .O(net_71845)
  );
  CEMux inmux_17_31_71851_71843 (
    .I(net_71851),
    .O(net_71843)
  );
  IoInMux inmux_17_31_71859_71837 (
    .I(net_71859),
    .O(net_71837)
  );
  ClkMux inmux_17_5_5_68715 (
    .I(net_5),
    .O(net_68715)
  );
  InMux inmux_17_5_68638_68671 (
    .I(net_68638),
    .O(net_68671)
  );
  InMux inmux_17_5_68645_68681 (
    .I(net_68645),
    .O(net_68681)
  );
  CEMux inmux_17_5_68646_68714 (
    .I(net_68646),
    .O(net_68714)
  );
  InMux inmux_17_5_68647_68705 (
    .I(net_68647),
    .O(net_68705)
  );
  InMux inmux_17_5_68648_68689 (
    .I(net_68648),
    .O(net_68689)
  );
  InMux inmux_17_5_68649_68712 (
    .I(net_68649),
    .O(net_68712)
  );
  InMux inmux_17_5_68650_68677 (
    .I(net_68650),
    .O(net_68677)
  );
  InMux inmux_17_5_68651_68670 (
    .I(net_68651),
    .O(net_68670)
  );
  InMux inmux_17_5_68651_68675 (
    .I(net_68651),
    .O(net_68675)
  );
  InMux inmux_17_5_68651_68680 (
    .I(net_68651),
    .O(net_68680)
  );
  InMux inmux_17_5_68651_68687 (
    .I(net_68651),
    .O(net_68687)
  );
  InMux inmux_17_5_68651_68706 (
    .I(net_68651),
    .O(net_68706)
  );
  InMux inmux_17_5_68651_68711 (
    .I(net_68651),
    .O(net_68711)
  );
  SRMux inmux_17_5_68655_68716 (
    .I(net_68655),
    .O(net_68716)
  );
  InMux inmux_17_5_68659_68698 (
    .I(net_68659),
    .O(net_68698)
  );
  InMux inmux_17_5_68662_68699 (
    .I(net_68662),
    .O(net_68699)
  );
  InMux inmux_17_5_68666_68701 (
    .I(net_68666),
    .O(net_68701)
  );
  ClkMux inmux_17_6_5_68838 (
    .I(net_5),
    .O(net_68838)
  );
  InMux inmux_17_6_68758_68834 (
    .I(net_68758),
    .O(net_68834)
  );
  InMux inmux_17_6_68759_68823 (
    .I(net_68759),
    .O(net_68823)
  );
  InMux inmux_17_6_68759_68833 (
    .I(net_68759),
    .O(net_68833)
  );
  InMux inmux_17_6_68764_68822 (
    .I(net_68764),
    .O(net_68822)
  );
  InMux inmux_17_6_68764_68836 (
    .I(net_68764),
    .O(net_68836)
  );
  InMux inmux_17_6_68766_68794 (
    .I(net_68766),
    .O(net_68794)
  );
  InMux inmux_17_6_68768_68816 (
    .I(net_68768),
    .O(net_68816)
  );
  InMux inmux_17_6_68768_68821 (
    .I(net_68768),
    .O(net_68821)
  );
  CEMux inmux_17_6_68769_68837 (
    .I(net_68769),
    .O(net_68837)
  );
  InMux inmux_17_6_68771_68815 (
    .I(net_68771),
    .O(net_68815)
  );
  InMux inmux_17_6_68773_68817 (
    .I(net_68773),
    .O(net_68817)
  );
  InMux inmux_17_6_68774_68824 (
    .I(net_68774),
    .O(net_68824)
  );
  InMux inmux_17_6_68781_68835 (
    .I(net_68781),
    .O(net_68835)
  );
  InMux inmux_17_6_68782_68792 (
    .I(net_68782),
    .O(net_68792)
  );
  SRMux inmux_17_6_68787_68839 (
    .I(net_68787),
    .O(net_68839)
  );
  ClkMux inmux_17_9_5_69207 (
    .I(net_5),
    .O(net_69207)
  );
  InMux inmux_17_9_69151_69166 (
    .I(net_69151),
    .O(net_69166)
  );
  CEMux inmux_17_9_8_69206 (
    .I(net_8),
    .O(net_69206)
  );
  ClkMux inmux_18_0_5_71874 (
    .I(net_5),
    .O(net_71874)
  );
  ClkMux inmux_18_0_5_71875 (
    .I(net_5),
    .O(net_71875)
  );
  CEMux inmux_18_0_71878_71873 (
    .I(net_71878),
    .O(net_71873)
  );
  IoInMux inmux_18_0_71885_71867 (
    .I(net_71885),
    .O(net_71867)
  );
  InMux inmux_18_10_73084_73132 (
    .I(net_73084),
    .O(net_73132)
  );
  InMux inmux_18_10_73085_73135 (
    .I(net_73085),
    .O(net_73135)
  );
  InMux inmux_18_10_73090_73133 (
    .I(net_73090),
    .O(net_73133)
  );
  InMux inmux_18_10_73105_73134 (
    .I(net_73105),
    .O(net_73134)
  );
  ClkMux inmux_18_12_5_73407 (
    .I(net_5),
    .O(net_73407)
  );
  InMux inmux_18_12_73330_73378 (
    .I(net_73330),
    .O(net_73378)
  );
  InMux inmux_18_12_73354_73396 (
    .I(net_73354),
    .O(net_73396)
  );
  InMux inmux_18_12_73355_73402 (
    .I(net_73355),
    .O(net_73402)
  );
  ClkMux inmux_18_13_5_73530 (
    .I(net_5),
    .O(net_73530)
  );
  InMux inmux_18_13_73452_73504 (
    .I(net_73452),
    .O(net_73504)
  );
  InMux inmux_18_13_73453_73503 (
    .I(net_73453),
    .O(net_73503)
  );
  InMux inmux_18_13_73454_73507 (
    .I(net_73454),
    .O(net_73507)
  );
  InMux inmux_18_13_73461_73492 (
    .I(net_73461),
    .O(net_73492)
  );
  InMux inmux_18_13_73462_73510 (
    .I(net_73462),
    .O(net_73510)
  );
  InMux inmux_18_13_73467_73527 (
    .I(net_73467),
    .O(net_73527)
  );
  InMux inmux_18_13_73473_73522 (
    .I(net_73473),
    .O(net_73522)
  );
  InMux inmux_18_13_73475_73502 (
    .I(net_73475),
    .O(net_73502)
  );
  InMux inmux_18_13_73475_73509 (
    .I(net_73475),
    .O(net_73509)
  );
  InMux inmux_18_13_73478_73484 (
    .I(net_73478),
    .O(net_73484)
  );
  InMux inmux_18_13_73479_73514 (
    .I(net_73479),
    .O(net_73514)
  );
  InMux inmux_18_13_73481_73497 (
    .I(net_73481),
    .O(net_73497)
  );
  CEMux inmux_18_14_10_73652 (
    .I(net_10),
    .O(net_73652)
  );
  SRMux inmux_18_14_11_73654 (
    .I(net_11),
    .O(net_73654)
  );
  ClkMux inmux_18_14_5_73653 (
    .I(net_5),
    .O(net_73653)
  );
  InMux inmux_18_14_73574_73607 (
    .I(net_73574),
    .O(net_73607)
  );
  InMux inmux_18_14_73575_73606 (
    .I(net_73575),
    .O(net_73606)
  );
  InMux inmux_18_14_73575_73613 (
    .I(net_73575),
    .O(net_73613)
  );
  InMux inmux_18_14_73575_73630 (
    .I(net_73575),
    .O(net_73630)
  );
  InMux inmux_18_14_73576_73633 (
    .I(net_73576),
    .O(net_73633)
  );
  InMux inmux_18_14_73580_73636 (
    .I(net_73580),
    .O(net_73636)
  );
  InMux inmux_18_14_73582_73608 (
    .I(net_73582),
    .O(net_73608)
  );
  InMux inmux_18_14_73583_73614 (
    .I(net_73583),
    .O(net_73614)
  );
  InMux inmux_18_14_73585_73650 (
    .I(net_73585),
    .O(net_73650)
  );
  InMux inmux_18_14_73588_73615 (
    .I(net_73588),
    .O(net_73615)
  );
  InMux inmux_18_14_73589_73625 (
    .I(net_73589),
    .O(net_73625)
  );
  InMux inmux_18_14_73590_73624 (
    .I(net_73590),
    .O(net_73624)
  );
  InMux inmux_18_14_73591_73618 (
    .I(net_73591),
    .O(net_73618)
  );
  InMux inmux_18_14_73591_73627 (
    .I(net_73591),
    .O(net_73627)
  );
  InMux inmux_18_14_73592_73619 (
    .I(net_73592),
    .O(net_73619)
  );
  InMux inmux_18_14_73595_73637 (
    .I(net_73595),
    .O(net_73637)
  );
  InMux inmux_18_14_73596_73621 (
    .I(net_73596),
    .O(net_73621)
  );
  InMux inmux_18_14_73599_73648 (
    .I(net_73599),
    .O(net_73648)
  );
  InMux inmux_18_14_73602_73632 (
    .I(net_73602),
    .O(net_73632)
  );
  InMux inmux_18_14_73604_73639 (
    .I(net_73604),
    .O(net_73639)
  );
  InMux inmux_18_14_73604_73651 (
    .I(net_73604),
    .O(net_73651)
  );
  ClkMux inmux_18_15_5_73776 (
    .I(net_5),
    .O(net_73776)
  );
  InMux inmux_18_15_73701_73732 (
    .I(net_73701),
    .O(net_73732)
  );
  InMux inmux_18_15_73713_73759 (
    .I(net_73713),
    .O(net_73759)
  );
  InMux inmux_18_15_73717_73744 (
    .I(net_73717),
    .O(net_73744)
  );
  InMux inmux_18_15_73722_73749 (
    .I(net_73722),
    .O(net_73749)
  );
  InMux inmux_18_15_73723_73767 (
    .I(net_73723),
    .O(net_73767)
  );
  InMux inmux_18_15_73724_73771 (
    .I(net_73724),
    .O(net_73771)
  );
  InMux inmux_18_15_73725_73753 (
    .I(net_73725),
    .O(net_73753)
  );
  ClkMux inmux_18_16_5_73899 (
    .I(net_5),
    .O(net_73899)
  );
  InMux inmux_18_16_73845_73867 (
    .I(net_73845),
    .O(net_73867)
  );
  InMux inmux_18_16_73849_73865 (
    .I(net_73849),
    .O(net_73865)
  );
  ClkMux inmux_18_17_5_74022 (
    .I(net_5),
    .O(net_74022)
  );
  InMux inmux_18_17_73946_74006 (
    .I(net_73946),
    .O(net_74006)
  );
  InMux inmux_18_17_73948_73987 (
    .I(net_73948),
    .O(net_73987)
  );
  InMux inmux_18_17_73950_74005 (
    .I(net_73950),
    .O(net_74005)
  );
  InMux inmux_18_17_73953_74013 (
    .I(net_73953),
    .O(net_74013)
  );
  InMux inmux_18_17_73955_74018 (
    .I(net_73955),
    .O(net_74018)
  );
  InMux inmux_18_17_73956_73978 (
    .I(net_73956),
    .O(net_73978)
  );
  InMux inmux_18_17_73962_74008 (
    .I(net_73962),
    .O(net_74008)
  );
  InMux inmux_18_17_73965_73983 (
    .I(net_73965),
    .O(net_73983)
  );
  InMux inmux_18_17_73969_74001 (
    .I(net_73969),
    .O(net_74001)
  );
  InMux inmux_18_17_73970_74007 (
    .I(net_73970),
    .O(net_74007)
  );
  InMux inmux_18_17_73971_73994 (
    .I(net_73971),
    .O(net_73994)
  );
  CEMux inmux_18_18_10_74144 (
    .I(net_10),
    .O(net_74144)
  );
  SRMux inmux_18_18_11_74146 (
    .I(net_11),
    .O(net_74146)
  );
  ClkMux inmux_18_18_5_74145 (
    .I(net_5),
    .O(net_74145)
  );
  InMux inmux_18_18_74065_74117 (
    .I(net_74065),
    .O(net_74117)
  );
  InMux inmux_18_18_74068_74125 (
    .I(net_74068),
    .O(net_74125)
  );
  InMux inmux_18_18_74070_74140 (
    .I(net_74070),
    .O(net_74140)
  );
  InMux inmux_18_18_74072_74113 (
    .I(net_74072),
    .O(net_74113)
  );
  InMux inmux_18_18_74074_74131 (
    .I(net_74074),
    .O(net_74131)
  );
  InMux inmux_18_18_74076_74112 (
    .I(net_74076),
    .O(net_74112)
  );
  InMux inmux_18_18_74076_74119 (
    .I(net_74076),
    .O(net_74119)
  );
  InMux inmux_18_18_74076_74129 (
    .I(net_74076),
    .O(net_74129)
  );
  InMux inmux_18_18_74076_74134 (
    .I(net_74076),
    .O(net_74134)
  );
  InMux inmux_18_18_74077_74135 (
    .I(net_74077),
    .O(net_74135)
  );
  InMux inmux_18_18_74080_74141 (
    .I(net_74080),
    .O(net_74141)
  );
  InMux inmux_18_18_74082_74116 (
    .I(net_74082),
    .O(net_74116)
  );
  InMux inmux_18_18_74083_74122 (
    .I(net_74083),
    .O(net_74122)
  );
  InMux inmux_18_18_74083_74143 (
    .I(net_74083),
    .O(net_74143)
  );
  InMux inmux_18_18_74084_74111 (
    .I(net_74084),
    .O(net_74111)
  );
  InMux inmux_18_18_74086_74128 (
    .I(net_74086),
    .O(net_74128)
  );
  InMux inmux_18_18_74091_74137 (
    .I(net_74091),
    .O(net_74137)
  );
  InMux inmux_18_18_74092_74124 (
    .I(net_74092),
    .O(net_74124)
  );
  CEMux inmux_18_19_10_74267 (
    .I(net_10),
    .O(net_74267)
  );
  ClkMux inmux_18_19_5_74268 (
    .I(net_5),
    .O(net_74268)
  );
  InMux inmux_18_19_74195_74263 (
    .I(net_74195),
    .O(net_74263)
  );
  ClkMux inmux_18_20_5_74391 (
    .I(net_5),
    .O(net_74391)
  );
  InMux inmux_18_20_74320_74387 (
    .I(net_74320),
    .O(net_74387)
  );
  ClkMux inmux_18_31_5_75675 (
    .I(net_5),
    .O(net_75675)
  );
  ClkMux inmux_18_31_5_75676 (
    .I(net_5),
    .O(net_75676)
  );
  CEMux inmux_18_31_75679_75674 (
    .I(net_75679),
    .O(net_75674)
  );
  IoInMux inmux_18_31_75682_75671 (
    .I(net_75682),
    .O(net_75671)
  );
  ClkMux inmux_18_5_5_72546 (
    .I(net_5),
    .O(net_72546)
  );
  InMux inmux_18_5_72466_72530 (
    .I(net_72466),
    .O(net_72530)
  );
  SRMux inmux_18_5_72479_72547 (
    .I(net_72479),
    .O(net_72547)
  );
  CEMux inmux_18_5_72484_72545 (
    .I(net_72484),
    .O(net_72545)
  );
  InMux inmux_18_5_72485_72541 (
    .I(net_72485),
    .O(net_72541)
  );
  InMux inmux_18_5_72495_72544 (
    .I(net_72495),
    .O(net_72544)
  );
  InMux inmux_18_5_72497_72532 (
    .I(net_72497),
    .O(net_72532)
  );
  ClkMux inmux_18_6_5_72669 (
    .I(net_5),
    .O(net_72669)
  );
  SRMux inmux_18_6_72593_72670 (
    .I(net_72593),
    .O(net_72670)
  );
  InMux inmux_18_6_72594_72635 (
    .I(net_72594),
    .O(net_72635)
  );
  InMux inmux_18_6_72594_72659 (
    .I(net_72594),
    .O(net_72659)
  );
  InMux inmux_18_6_72596_72652 (
    .I(net_72596),
    .O(net_72652)
  );
  InMux inmux_18_6_72597_72664 (
    .I(net_72597),
    .O(net_72664)
  );
  CEMux inmux_18_6_72600_72668 (
    .I(net_72600),
    .O(net_72668)
  );
  InMux inmux_18_6_72601_72630 (
    .I(net_72601),
    .O(net_72630)
  );
  InMux inmux_18_6_72602_72624 (
    .I(net_72602),
    .O(net_72624)
  );
  InMux inmux_18_6_72602_72653 (
    .I(net_72602),
    .O(net_72653)
  );
  InMux inmux_18_6_72604_72629 (
    .I(net_72604),
    .O(net_72629)
  );
  InMux inmux_18_6_72605_72631 (
    .I(net_72605),
    .O(net_72631)
  );
  InMux inmux_18_6_72607_72622 (
    .I(net_72607),
    .O(net_72622)
  );
  InMux inmux_18_6_72607_72655 (
    .I(net_72607),
    .O(net_72655)
  );
  InMux inmux_18_6_72610_72625 (
    .I(net_72610),
    .O(net_72625)
  );
  InMux inmux_18_6_72610_72628 (
    .I(net_72610),
    .O(net_72628)
  );
  InMux inmux_18_6_72610_72654 (
    .I(net_72610),
    .O(net_72654)
  );
  InMux inmux_18_6_72612_72637 (
    .I(net_72612),
    .O(net_72637)
  );
  InMux inmux_18_6_72612_72666 (
    .I(net_72612),
    .O(net_72666)
  );
  InMux inmux_18_6_72613_72661 (
    .I(net_72613),
    .O(net_72661)
  );
  InMux inmux_18_6_72618_72660 (
    .I(net_72618),
    .O(net_72660)
  );
  ClkMux inmux_19_13_5_77086 (
    .I(net_5),
    .O(net_77086)
  );
  InMux inmux_19_13_77027_77091 (
    .I(net_77027),
    .O(net_77091)
  );
  InMux inmux_19_13_77030_77078 (
    .I(net_77030),
    .O(net_77078)
  );
  InMux inmux_19_13_77031_77095 (
    .I(net_77031),
    .O(net_77095)
  );
  InMux inmux_19_13_77033_77089 (
    .I(net_77033),
    .O(net_77089)
  );
  InMux inmux_19_13_77034_77080 (
    .I(net_77034),
    .O(net_77080)
  );
  InMux inmux_19_13_77035_77096 (
    .I(net_77035),
    .O(net_77096)
  );
  InMux inmux_19_13_77036_77076 (
    .I(net_77036),
    .O(net_77076)
  );
  InMux inmux_19_13_77038_77079 (
    .I(net_77038),
    .O(net_77079)
  );
  InMux inmux_19_13_77039_77092 (
    .I(net_77039),
    .O(net_77092)
  );
  InMux inmux_19_13_77040_77081 (
    .I(net_77040),
    .O(net_77081)
  );
  InMux inmux_19_13_77042_77083 (
    .I(net_77042),
    .O(net_77083)
  );
  InMux inmux_19_13_77044_77090 (
    .I(net_77044),
    .O(net_77090)
  );
  InMux inmux_19_13_77048_77075 (
    .I(net_77048),
    .O(net_77075)
  );
  InMux inmux_19_13_77049_77093 (
    .I(net_77049),
    .O(net_77093)
  );
  InMux inmux_19_13_77050_77094 (
    .I(net_77050),
    .O(net_77094)
  );
  CEMux inmux_19_13_77054_77087 (
    .I(net_77054),
    .O(net_77087)
  );
  SRMux inmux_19_13_77056_77088 (
    .I(net_77056),
    .O(net_77088)
  );
  InMux inmux_19_13_77057_77082 (
    .I(net_77057),
    .O(net_77082)
  );
  ClkMux inmux_19_14_5_77188 (
    .I(net_5),
    .O(net_77188)
  );
  InMux inmux_19_14_77129_77190 (
    .I(net_77129),
    .O(net_77190)
  );
  InMux inmux_19_14_77130_77193 (
    .I(net_77130),
    .O(net_77193)
  );
  InMux inmux_19_14_77131_77178 (
    .I(net_77131),
    .O(net_77178)
  );
  InMux inmux_19_14_77132_77182 (
    .I(net_77132),
    .O(net_77182)
  );
  InMux inmux_19_14_77133_77192 (
    .I(net_77133),
    .O(net_77192)
  );
  InMux inmux_19_14_77134_77197 (
    .I(net_77134),
    .O(net_77197)
  );
  InMux inmux_19_14_77135_77181 (
    .I(net_77135),
    .O(net_77181)
  );
  InMux inmux_19_14_77137_77184 (
    .I(net_77137),
    .O(net_77184)
  );
  InMux inmux_19_14_77141_77191 (
    .I(net_77141),
    .O(net_77191)
  );
  SRMux inmux_19_14_77142_77198 (
    .I(net_77142),
    .O(net_77198)
  );
  InMux inmux_19_14_77147_77183 (
    .I(net_77147),
    .O(net_77183)
  );
  InMux inmux_19_14_77150_77177 (
    .I(net_77150),
    .O(net_77177)
  );
  InMux inmux_19_14_77151_77185 (
    .I(net_77151),
    .O(net_77185)
  );
  InMux inmux_19_14_77152_77195 (
    .I(net_77152),
    .O(net_77195)
  );
  CEMux inmux_19_14_77156_77189 (
    .I(net_77156),
    .O(net_77189)
  );
  InMux inmux_19_14_77157_77180 (
    .I(net_77157),
    .O(net_77180)
  );
  InMux inmux_19_14_77158_77194 (
    .I(net_77158),
    .O(net_77194)
  );
  InMux inmux_19_14_77160_77196 (
    .I(net_77160),
    .O(net_77196)
  );
  ClkMux inmux_19_15_5_77290 (
    .I(net_5),
    .O(net_77290)
  );
  InMux inmux_19_15_77231_77297 (
    .I(net_77231),
    .O(net_77297)
  );
  InMux inmux_19_15_77232_77286 (
    .I(net_77232),
    .O(net_77286)
  );
  CEMux inmux_19_15_77233_77291 (
    .I(net_77233),
    .O(net_77291)
  );
  InMux inmux_19_15_77234_77296 (
    .I(net_77234),
    .O(net_77296)
  );
  SRMux inmux_19_15_77235_77292 (
    .I(net_77235),
    .O(net_77292)
  );
  InMux inmux_19_15_77236_77279 (
    .I(net_77236),
    .O(net_77279)
  );
  InMux inmux_19_15_77239_77294 (
    .I(net_77239),
    .O(net_77294)
  );
  InMux inmux_19_15_77240_77299 (
    .I(net_77240),
    .O(net_77299)
  );
  InMux inmux_19_15_77246_77280 (
    .I(net_77246),
    .O(net_77280)
  );
  InMux inmux_19_15_77247_77283 (
    .I(net_77247),
    .O(net_77283)
  );
  InMux inmux_19_15_77248_77282 (
    .I(net_77248),
    .O(net_77282)
  );
  InMux inmux_19_15_77251_77287 (
    .I(net_77251),
    .O(net_77287)
  );
  InMux inmux_19_15_77252_77284 (
    .I(net_77252),
    .O(net_77284)
  );
  InMux inmux_19_15_77254_77300 (
    .I(net_77254),
    .O(net_77300)
  );
  InMux inmux_19_15_77258_77293 (
    .I(net_77258),
    .O(net_77293)
  );
  InMux inmux_19_15_77260_77295 (
    .I(net_77260),
    .O(net_77295)
  );
  InMux inmux_19_15_77261_77298 (
    .I(net_77261),
    .O(net_77298)
  );
  InMux inmux_19_15_77262_77285 (
    .I(net_77262),
    .O(net_77285)
  );
  ClkMux inmux_19_16_5_77392 (
    .I(net_5),
    .O(net_77392)
  );
  InMux inmux_19_16_77334_77395 (
    .I(net_77334),
    .O(net_77395)
  );
  InMux inmux_19_16_77339_77394 (
    .I(net_77339),
    .O(net_77394)
  );
  InMux inmux_19_16_77342_77396 (
    .I(net_77342),
    .O(net_77396)
  );
  InMux inmux_19_16_77343_77381 (
    .I(net_77343),
    .O(net_77381)
  );
  InMux inmux_19_16_77346_77398 (
    .I(net_77346),
    .O(net_77398)
  );
  InMux inmux_19_16_77349_77400 (
    .I(net_77349),
    .O(net_77400)
  );
  CEMux inmux_19_16_77351_77393 (
    .I(net_77351),
    .O(net_77393)
  );
  SRMux inmux_19_16_77353_77402 (
    .I(net_77353),
    .O(net_77402)
  );
  InMux inmux_19_16_77354_77399 (
    .I(net_77354),
    .O(net_77399)
  );
  InMux inmux_19_16_77356_77401 (
    .I(net_77356),
    .O(net_77401)
  );
  InMux inmux_19_16_77357_77397 (
    .I(net_77357),
    .O(net_77397)
  );
  InMux inmux_19_16_77358_77382 (
    .I(net_77358),
    .O(net_77382)
  );
  InMux inmux_19_16_77359_77384 (
    .I(net_77359),
    .O(net_77384)
  );
  InMux inmux_19_16_77360_77385 (
    .I(net_77360),
    .O(net_77385)
  );
  InMux inmux_19_16_77361_77386 (
    .I(net_77361),
    .O(net_77386)
  );
  InMux inmux_19_16_77362_77387 (
    .I(net_77362),
    .O(net_77387)
  );
  InMux inmux_19_16_77363_77388 (
    .I(net_77363),
    .O(net_77388)
  );
  InMux inmux_19_16_77364_77389 (
    .I(net_77364),
    .O(net_77389)
  );
  ClkMux inmux_19_17_5_77494 (
    .I(net_5),
    .O(net_77494)
  );
  InMux inmux_19_17_77435_77503 (
    .I(net_77435),
    .O(net_77503)
  );
  InMux inmux_19_17_77436_77486 (
    .I(net_77436),
    .O(net_77486)
  );
  InMux inmux_19_17_77437_77484 (
    .I(net_77437),
    .O(net_77484)
  );
  InMux inmux_19_17_77439_77497 (
    .I(net_77439),
    .O(net_77497)
  );
  InMux inmux_19_17_77440_77488 (
    .I(net_77440),
    .O(net_77488)
  );
  InMux inmux_19_17_77446_77487 (
    .I(net_77446),
    .O(net_77487)
  );
  InMux inmux_19_17_77447_77504 (
    .I(net_77447),
    .O(net_77504)
  );
  InMux inmux_19_17_77449_77498 (
    .I(net_77449),
    .O(net_77498)
  );
  InMux inmux_19_17_77450_77489 (
    .I(net_77450),
    .O(net_77489)
  );
  InMux inmux_19_17_77452_77490 (
    .I(net_77452),
    .O(net_77490)
  );
  InMux inmux_19_17_77453_77501 (
    .I(net_77453),
    .O(net_77501)
  );
  InMux inmux_19_17_77456_77483 (
    .I(net_77456),
    .O(net_77483)
  );
  InMux inmux_19_17_77457_77491 (
    .I(net_77457),
    .O(net_77491)
  );
  InMux inmux_19_17_77461_77500 (
    .I(net_77461),
    .O(net_77500)
  );
  CEMux inmux_19_17_77462_77495 (
    .I(net_77462),
    .O(net_77495)
  );
  SRMux inmux_19_17_77464_77496 (
    .I(net_77464),
    .O(net_77496)
  );
  InMux inmux_19_17_77466_77499 (
    .I(net_77466),
    .O(net_77499)
  );
  ClkMux inmux_19_18_5_77596 (
    .I(net_5),
    .O(net_77596)
  );
  InMux inmux_19_18_77538_77588 (
    .I(net_77538),
    .O(net_77588)
  );
  CEMux inmux_19_18_77539_77597 (
    .I(net_77539),
    .O(net_77597)
  );
  InMux inmux_19_18_77541_77600 (
    .I(net_77541),
    .O(net_77600)
  );
  InMux inmux_19_18_77542_77585 (
    .I(net_77542),
    .O(net_77585)
  );
  InMux inmux_19_18_77545_77605 (
    .I(net_77545),
    .O(net_77605)
  );
  InMux inmux_19_18_77548_77602 (
    .I(net_77548),
    .O(net_77602)
  );
  InMux inmux_19_18_77549_77592 (
    .I(net_77549),
    .O(net_77592)
  );
  SRMux inmux_19_18_77550_77606 (
    .I(net_77550),
    .O(net_77606)
  );
  InMux inmux_19_18_77553_77591 (
    .I(net_77553),
    .O(net_77591)
  );
  InMux inmux_19_18_77555_77586 (
    .I(net_77555),
    .O(net_77586)
  );
  InMux inmux_19_18_77558_77599 (
    .I(net_77558),
    .O(net_77599)
  );
  InMux inmux_19_18_77559_77589 (
    .I(net_77559),
    .O(net_77589)
  );
  InMux inmux_19_18_77561_77590 (
    .I(net_77561),
    .O(net_77590)
  );
  InMux inmux_19_18_77562_77598 (
    .I(net_77562),
    .O(net_77598)
  );
  InMux inmux_19_18_77563_77603 (
    .I(net_77563),
    .O(net_77603)
  );
  InMux inmux_19_18_77564_77604 (
    .I(net_77564),
    .O(net_77604)
  );
  InMux inmux_19_18_77565_77601 (
    .I(net_77565),
    .O(net_77601)
  );
  InMux inmux_19_18_77568_77593 (
    .I(net_77568),
    .O(net_77593)
  );
  InMux inmux_1_30_11035_11052 (
    .I(net_11035),
    .O(net_11052)
  );
  ClkMux inmux_20_10_5_80192 (
    .I(net_5),
    .O(net_80192)
  );
  CEMux inmux_20_10_80114_80191 (
    .I(net_80114),
    .O(net_80191)
  );
  InMux inmux_20_10_80117_80177 (
    .I(net_80117),
    .O(net_80177)
  );
  InMux inmux_20_10_80117_80189 (
    .I(net_80117),
    .O(net_80189)
  );
  InMux inmux_20_10_80119_80148 (
    .I(net_80119),
    .O(net_80148)
  );
  InMux inmux_20_10_80119_80187 (
    .I(net_80119),
    .O(net_80187)
  );
  InMux inmux_20_10_80121_80164 (
    .I(net_80121),
    .O(net_80164)
  );
  InMux inmux_20_10_80122_80165 (
    .I(net_80122),
    .O(net_80165)
  );
  InMux inmux_20_10_80123_80178 (
    .I(net_80123),
    .O(net_80178)
  );
  SRMux inmux_20_10_80125_80193 (
    .I(net_80125),
    .O(net_80193)
  );
  InMux inmux_20_10_80129_80163 (
    .I(net_80129),
    .O(net_80163)
  );
  InMux inmux_20_10_80132_80176 (
    .I(net_80132),
    .O(net_80176)
  );
  InMux inmux_20_10_80136_80175 (
    .I(net_80136),
    .O(net_80175)
  );
  InMux inmux_20_10_80137_80147 (
    .I(net_80137),
    .O(net_80147)
  );
  InMux inmux_20_10_80139_80166 (
    .I(net_80139),
    .O(net_80166)
  );
  InMux inmux_20_10_80140_80146 (
    .I(net_80140),
    .O(net_80146)
  );
  ClkMux inmux_20_11_5_80315 (
    .I(net_5),
    .O(net_80315)
  );
  InMux inmux_20_11_80242_80300 (
    .I(net_80242),
    .O(net_80300)
  );
  CEMux inmux_20_12_10_80437 (
    .I(net_10),
    .O(net_80437)
  );
  SRMux inmux_20_12_11_80439 (
    .I(net_11),
    .O(net_80439)
  );
  ClkMux inmux_20_12_5_80438 (
    .I(net_5),
    .O(net_80438)
  );
  InMux inmux_20_12_80359_80397 (
    .I(net_80359),
    .O(net_80397)
  );
  InMux inmux_20_12_80359_80404 (
    .I(net_80359),
    .O(net_80404)
  );
  InMux inmux_20_12_80359_80409 (
    .I(net_80359),
    .O(net_80409)
  );
  InMux inmux_20_12_80359_80421 (
    .I(net_80359),
    .O(net_80421)
  );
  InMux inmux_20_12_80359_80428 (
    .I(net_80359),
    .O(net_80428)
  );
  InMux inmux_20_12_80360_80424 (
    .I(net_80360),
    .O(net_80424)
  );
  InMux inmux_20_12_80364_80400 (
    .I(net_80364),
    .O(net_80400)
  );
  InMux inmux_20_12_80368_80435 (
    .I(net_80368),
    .O(net_80435)
  );
  InMux inmux_20_12_80369_80415 (
    .I(net_80369),
    .O(net_80415)
  );
  InMux inmux_20_12_80371_80405 (
    .I(net_80371),
    .O(net_80405)
  );
  InMux inmux_20_12_80372_80392 (
    .I(net_80372),
    .O(net_80392)
  );
  InMux inmux_20_12_80373_80422 (
    .I(net_80373),
    .O(net_80422)
  );
  InMux inmux_20_12_80375_80433 (
    .I(net_80375),
    .O(net_80433)
  );
  InMux inmux_20_12_80376_80393 (
    .I(net_80376),
    .O(net_80393)
  );
  InMux inmux_20_12_80376_80417 (
    .I(net_80376),
    .O(net_80417)
  );
  InMux inmux_20_12_80376_80436 (
    .I(net_80376),
    .O(net_80436)
  );
  InMux inmux_20_12_80377_80430 (
    .I(net_80377),
    .O(net_80430)
  );
  InMux inmux_20_12_80378_80429 (
    .I(net_80378),
    .O(net_80429)
  );
  InMux inmux_20_12_80379_80418 (
    .I(net_80379),
    .O(net_80418)
  );
  InMux inmux_20_12_80380_80398 (
    .I(net_80380),
    .O(net_80398)
  );
  InMux inmux_20_12_80381_80406 (
    .I(net_80381),
    .O(net_80406)
  );
  InMux inmux_20_12_80385_80412 (
    .I(net_80385),
    .O(net_80412)
  );
  InMux inmux_20_12_80388_80394 (
    .I(net_80388),
    .O(net_80394)
  );
  InMux inmux_20_12_80389_80410 (
    .I(net_80389),
    .O(net_80410)
  );
  CEMux inmux_20_13_10_80560 (
    .I(net_10),
    .O(net_80560)
  );
  SRMux inmux_20_13_11_80562 (
    .I(net_11),
    .O(net_80562)
  );
  ClkMux inmux_20_13_5_80561 (
    .I(net_5),
    .O(net_80561)
  );
  InMux inmux_20_13_80481_80552 (
    .I(net_80481),
    .O(net_80552)
  );
  InMux inmux_20_13_80482_80539 (
    .I(net_80482),
    .O(net_80539)
  );
  InMux inmux_20_13_80483_80523 (
    .I(net_80483),
    .O(net_80523)
  );
  InMux inmux_20_13_80485_80528 (
    .I(net_80485),
    .O(net_80528)
  );
  InMux inmux_20_13_80486_80529 (
    .I(net_80486),
    .O(net_80529)
  );
  InMux inmux_20_13_80489_80544 (
    .I(net_80489),
    .O(net_80544)
  );
  InMux inmux_20_13_80491_80532 (
    .I(net_80491),
    .O(net_80532)
  );
  InMux inmux_20_13_80492_80516 (
    .I(net_80492),
    .O(net_80516)
  );
  InMux inmux_20_13_80493_80515 (
    .I(net_80493),
    .O(net_80515)
  );
  InMux inmux_20_13_80494_80514 (
    .I(net_80494),
    .O(net_80514)
  );
  InMux inmux_20_13_80495_80517 (
    .I(net_80495),
    .O(net_80517)
  );
  InMux inmux_20_13_80499_80545 (
    .I(net_80499),
    .O(net_80545)
  );
  InMux inmux_20_13_80501_80521 (
    .I(net_80501),
    .O(net_80521)
  );
  InMux inmux_20_13_80501_80526 (
    .I(net_80501),
    .O(net_80526)
  );
  InMux inmux_20_13_80501_80533 (
    .I(net_80501),
    .O(net_80533)
  );
  InMux inmux_20_13_80501_80540 (
    .I(net_80501),
    .O(net_80540)
  );
  InMux inmux_20_13_80501_80547 (
    .I(net_80501),
    .O(net_80547)
  );
  InMux inmux_20_13_80501_80550 (
    .I(net_80501),
    .O(net_80550)
  );
  InMux inmux_20_13_80501_80557 (
    .I(net_80501),
    .O(net_80557)
  );
  InMux inmux_20_13_80502_80522 (
    .I(net_80502),
    .O(net_80522)
  );
  InMux inmux_20_13_80503_80535 (
    .I(net_80503),
    .O(net_80535)
  );
  InMux inmux_20_13_80507_80556 (
    .I(net_80507),
    .O(net_80556)
  );
  InMux inmux_20_13_80509_80558 (
    .I(net_80509),
    .O(net_80558)
  );
  InMux inmux_20_13_80510_80538 (
    .I(net_80510),
    .O(net_80538)
  );
  InMux inmux_20_13_80511_80551 (
    .I(net_80511),
    .O(net_80551)
  );
  ClkMux inmux_20_14_5_80684 (
    .I(net_5),
    .O(net_80684)
  );
  InMux inmux_20_14_80604_80656 (
    .I(net_80604),
    .O(net_80656)
  );
  InMux inmux_20_14_80604_80680 (
    .I(net_80604),
    .O(net_80680)
  );
  InMux inmux_20_14_80605_80638 (
    .I(net_80605),
    .O(net_80638)
  );
  InMux inmux_20_14_80605_80669 (
    .I(net_80605),
    .O(net_80669)
  );
  InMux inmux_20_14_80605_80674 (
    .I(net_80605),
    .O(net_80674)
  );
  InMux inmux_20_14_80609_80681 (
    .I(net_80609),
    .O(net_80681)
  );
  InMux inmux_20_14_80611_80667 (
    .I(net_80611),
    .O(net_80667)
  );
  InMux inmux_20_14_80612_80657 (
    .I(net_80612),
    .O(net_80657)
  );
  InMux inmux_20_14_80613_80639 (
    .I(net_80613),
    .O(net_80639)
  );
  InMux inmux_20_14_80618_80664 (
    .I(net_80618),
    .O(net_80664)
  );
  InMux inmux_20_14_80619_80637 (
    .I(net_80619),
    .O(net_80637)
  );
  InMux inmux_20_14_80620_80673 (
    .I(net_80620),
    .O(net_80673)
  );
  InMux inmux_20_14_80622_80670 (
    .I(net_80622),
    .O(net_80670)
  );
  InMux inmux_20_14_80623_80676 (
    .I(net_80623),
    .O(net_80676)
  );
  InMux inmux_20_14_80624_80658 (
    .I(net_80624),
    .O(net_80658)
  );
  InMux inmux_20_14_80626_80682 (
    .I(net_80626),
    .O(net_80682)
  );
  InMux inmux_20_14_80628_80655 (
    .I(net_80628),
    .O(net_80655)
  );
  InMux inmux_20_14_80628_80679 (
    .I(net_80628),
    .O(net_80679)
  );
  InMux inmux_20_14_80631_80649 (
    .I(net_80631),
    .O(net_80649)
  );
  InMux inmux_20_14_80635_80644 (
    .I(net_80635),
    .O(net_80644)
  );
  CEMux inmux_20_15_10_80806 (
    .I(net_10),
    .O(net_80806)
  );
  SRMux inmux_20_15_11_80808 (
    .I(net_11),
    .O(net_80808)
  );
  ClkMux inmux_20_15_5_80807 (
    .I(net_5),
    .O(net_80807)
  );
  InMux inmux_20_15_80727_80779 (
    .I(net_80727),
    .O(net_80779)
  );
  InMux inmux_20_15_80729_80774 (
    .I(net_80729),
    .O(net_80774)
  );
  InMux inmux_20_15_80731_80760 (
    .I(net_80731),
    .O(net_80760)
  );
  InMux inmux_20_15_80735_80778 (
    .I(net_80735),
    .O(net_80778)
  );
  InMux inmux_20_15_80736_80805 (
    .I(net_80736),
    .O(net_80805)
  );
  InMux inmux_20_15_80738_80798 (
    .I(net_80738),
    .O(net_80798)
  );
  InMux inmux_20_15_80739_80761 (
    .I(net_80739),
    .O(net_80761)
  );
  InMux inmux_20_15_80740_80784 (
    .I(net_80740),
    .O(net_80784)
  );
  InMux inmux_20_15_80741_80804 (
    .I(net_80741),
    .O(net_80804)
  );
  InMux inmux_20_15_80743_80772 (
    .I(net_80743),
    .O(net_80772)
  );
  InMux inmux_20_15_80744_80775 (
    .I(net_80744),
    .O(net_80775)
  );
  InMux inmux_20_15_80744_80780 (
    .I(net_80744),
    .O(net_80780)
  );
  InMux inmux_20_15_80744_80787 (
    .I(net_80744),
    .O(net_80787)
  );
  InMux inmux_20_15_80744_80799 (
    .I(net_80744),
    .O(net_80799)
  );
  InMux inmux_20_15_80744_80802 (
    .I(net_80744),
    .O(net_80802)
  );
  InMux inmux_20_15_80745_80762 (
    .I(net_80745),
    .O(net_80762)
  );
  InMux inmux_20_15_80747_80767 (
    .I(net_80747),
    .O(net_80767)
  );
  InMux inmux_20_15_80749_80791 (
    .I(net_80749),
    .O(net_80791)
  );
  InMux inmux_20_15_80751_80797 (
    .I(net_80751),
    .O(net_80797)
  );
  InMux inmux_20_15_80752_80769 (
    .I(net_80752),
    .O(net_80769)
  );
  InMux inmux_20_15_80752_80793 (
    .I(net_80752),
    .O(net_80793)
  );
  InMux inmux_20_15_80753_80768 (
    .I(net_80753),
    .O(net_80768)
  );
  InMux inmux_20_15_80755_80790 (
    .I(net_80755),
    .O(net_80790)
  );
  InMux inmux_20_15_80757_80785 (
    .I(net_80757),
    .O(net_80785)
  );
  ClkMux inmux_20_16_5_80930 (
    .I(net_5),
    .O(net_80930)
  );
  InMux inmux_20_16_80855_80884 (
    .I(net_80855),
    .O(net_80884)
  );
  InMux inmux_20_16_80859_80890 (
    .I(net_80859),
    .O(net_80890)
  );
  InMux inmux_20_16_80862_80908 (
    .I(net_80862),
    .O(net_80908)
  );
  InMux inmux_20_16_80864_80920 (
    .I(net_80864),
    .O(net_80920)
  );
  InMux inmux_20_16_80868_80897 (
    .I(net_80868),
    .O(net_80897)
  );
  InMux inmux_20_16_80870_80885 (
    .I(net_80870),
    .O(net_80885)
  );
  InMux inmux_20_16_80871_80915 (
    .I(net_80871),
    .O(net_80915)
  );
  InMux inmux_20_16_80877_80902 (
    .I(net_80877),
    .O(net_80902)
  );
  InMux inmux_20_16_80881_80926 (
    .I(net_80881),
    .O(net_80926)
  );
  InMux inmux_20_16_80882_80892 (
    .I(net_80882),
    .O(net_80892)
  );
  InMux inmux_20_16_80888_80898 (
    .I(net_80888),
    .O(net_80898)
  );
  InMux inmux_20_16_80894_80904 (
    .I(net_80894),
    .O(net_80904)
  );
  InMux inmux_20_16_80900_80910 (
    .I(net_80900),
    .O(net_80910)
  );
  InMux inmux_20_16_80906_80916 (
    .I(net_80906),
    .O(net_80916)
  );
  InMux inmux_20_16_80912_80922 (
    .I(net_80912),
    .O(net_80922)
  );
  InMux inmux_20_16_80918_80928 (
    .I(net_80918),
    .O(net_80928)
  );
  CEMux inmux_20_17_10_81052 (
    .I(net_10),
    .O(net_81052)
  );
  SRMux inmux_20_17_11_81054 (
    .I(net_11),
    .O(net_81054)
  );
  ClkMux inmux_20_17_5_81053 (
    .I(net_5),
    .O(net_81053)
  );
  InMux inmux_20_17_80975_81025 (
    .I(net_80975),
    .O(net_81025)
  );
  InMux inmux_20_17_80976_81036 (
    .I(net_80976),
    .O(net_81036)
  );
  InMux inmux_20_17_80977_81018 (
    .I(net_80977),
    .O(net_81018)
  );
  InMux inmux_20_17_80978_81019 (
    .I(net_80978),
    .O(net_81019)
  );
  InMux inmux_20_17_80979_81008 (
    .I(net_80979),
    .O(net_81008)
  );
  InMux inmux_20_17_80980_81033 (
    .I(net_80980),
    .O(net_81033)
  );
  InMux inmux_20_17_80984_81030 (
    .I(net_80984),
    .O(net_81030)
  );
  InMux inmux_20_17_80985_81050 (
    .I(net_80985),
    .O(net_81050)
  );
  InMux inmux_20_17_80986_81006 (
    .I(net_80986),
    .O(net_81006)
  );
  InMux inmux_20_17_80986_81032 (
    .I(net_80986),
    .O(net_81032)
  );
  InMux inmux_20_17_80987_81045 (
    .I(net_80987),
    .O(net_81045)
  );
  InMux inmux_20_17_80989_81015 (
    .I(net_80989),
    .O(net_81015)
  );
  InMux inmux_20_17_80990_81007 (
    .I(net_80990),
    .O(net_81007)
  );
  InMux inmux_20_17_80990_81031 (
    .I(net_80990),
    .O(net_81031)
  );
  InMux inmux_20_17_80991_81051 (
    .I(net_80991),
    .O(net_81051)
  );
  InMux inmux_20_17_80992_81009 (
    .I(net_80992),
    .O(net_81009)
  );
  InMux inmux_20_17_80993_81020 (
    .I(net_80993),
    .O(net_81020)
  );
  InMux inmux_20_17_80995_81039 (
    .I(net_80995),
    .O(net_81039)
  );
  InMux inmux_20_17_80996_81043 (
    .I(net_80996),
    .O(net_81043)
  );
  InMux inmux_20_17_80997_81012 (
    .I(net_80997),
    .O(net_81012)
  );
  InMux inmux_20_17_80998_81027 (
    .I(net_80998),
    .O(net_81027)
  );
  InMux inmux_20_17_81001_81021 (
    .I(net_81001),
    .O(net_81021)
  );
  InMux inmux_20_17_81002_81044 (
    .I(net_81002),
    .O(net_81044)
  );
  InMux inmux_20_17_81003_81014 (
    .I(net_81003),
    .O(net_81014)
  );
  InMux inmux_20_17_81003_81024 (
    .I(net_81003),
    .O(net_81024)
  );
  InMux inmux_20_17_81003_81038 (
    .I(net_81003),
    .O(net_81038)
  );
  InMux inmux_20_17_81003_81048 (
    .I(net_81003),
    .O(net_81048)
  );
  CEMux inmux_20_18_10_81175 (
    .I(net_10),
    .O(net_81175)
  );
  SRMux inmux_20_18_11_81177 (
    .I(net_11),
    .O(net_81177)
  );
  ClkMux inmux_20_18_5_81176 (
    .I(net_5),
    .O(net_81176)
  );
  InMux inmux_20_18_81098_81150 (
    .I(net_81098),
    .O(net_81150)
  );
  InMux inmux_20_18_81099_81135 (
    .I(net_81099),
    .O(net_81135)
  );
  InMux inmux_20_18_81102_81138 (
    .I(net_81102),
    .O(net_81138)
  );
  InMux inmux_20_18_81102_81148 (
    .I(net_81102),
    .O(net_81148)
  );
  InMux inmux_20_18_81102_81153 (
    .I(net_81102),
    .O(net_81153)
  );
  InMux inmux_20_18_81102_81174 (
    .I(net_81102),
    .O(net_81174)
  );
  InMux inmux_20_18_81103_81154 (
    .I(net_81103),
    .O(net_81154)
  );
  InMux inmux_20_18_81105_81162 (
    .I(net_81105),
    .O(net_81162)
  );
  InMux inmux_20_18_81107_81155 (
    .I(net_81107),
    .O(net_81155)
  );
  InMux inmux_20_18_81110_81173 (
    .I(net_81110),
    .O(net_81173)
  );
  InMux inmux_20_18_81111_81136 (
    .I(net_81111),
    .O(net_81136)
  );
  InMux inmux_20_18_81112_81160 (
    .I(net_81112),
    .O(net_81160)
  );
  InMux inmux_20_18_81115_81149 (
    .I(net_81115),
    .O(net_81149)
  );
  InMux inmux_20_18_81119_81161 (
    .I(net_81119),
    .O(net_81161)
  );
  InMux inmux_20_18_81120_81159 (
    .I(net_81120),
    .O(net_81159)
  );
  InMux inmux_20_18_81125_81172 (
    .I(net_81125),
    .O(net_81172)
  );
  ClkMux inmux_20_19_5_81299 (
    .I(net_5),
    .O(net_81299)
  );
  InMux inmux_20_19_81236_81289 (
    .I(net_81236),
    .O(net_81289)
  );
  InMux inmux_20_19_81240_81294 (
    .I(net_81240),
    .O(net_81294)
  );
  ClkMux inmux_20_6_5_79700 (
    .I(net_5),
    .O(net_79700)
  );
  CEMux inmux_20_6_79622_79699 (
    .I(net_79622),
    .O(net_79699)
  );
  InMux inmux_20_6_79624_79655 (
    .I(net_79624),
    .O(net_79655)
  );
  InMux inmux_20_6_79628_79656 (
    .I(net_79628),
    .O(net_79656)
  );
  InMux inmux_20_6_79630_79697 (
    .I(net_79630),
    .O(net_79697)
  );
  InMux inmux_20_6_79635_79667 (
    .I(net_79635),
    .O(net_79667)
  );
  InMux inmux_20_6_79635_79686 (
    .I(net_79635),
    .O(net_79686)
  );
  InMux inmux_20_6_79638_79653 (
    .I(net_79638),
    .O(net_79653)
  );
  InMux inmux_20_6_79641_79668 (
    .I(net_79641),
    .O(net_79668)
  );
  InMux inmux_20_6_79641_79685 (
    .I(net_79641),
    .O(net_79685)
  );
  InMux inmux_20_6_79646_79654 (
    .I(net_79646),
    .O(net_79654)
  );
  SRMux inmux_20_6_79649_79701 (
    .I(net_79649),
    .O(net_79701)
  );
  InMux inmux_20_7_79756_79778 (
    .I(net_79756),
    .O(net_79778)
  );
  InMux inmux_20_7_79761_79776 (
    .I(net_79761),
    .O(net_79776)
  );
  ClkMux inmux_20_9_5_80069 (
    .I(net_5),
    .O(net_80069)
  );
  CEMux inmux_20_9_79991_80068 (
    .I(net_79991),
    .O(net_80068)
  );
  InMux inmux_20_9_79997_80025 (
    .I(net_79997),
    .O(net_80025)
  );
  InMux inmux_20_9_79997_80028 (
    .I(net_79997),
    .O(net_80028)
  );
  InMux inmux_20_9_80000_80022 (
    .I(net_80000),
    .O(net_80022)
  );
  InMux inmux_20_9_80004_80053 (
    .I(net_80004),
    .O(net_80053)
  );
  InMux inmux_20_9_80014_80055 (
    .I(net_80014),
    .O(net_80055)
  );
  ClkMux inmux_21_10_5_84023 (
    .I(net_5),
    .O(net_84023)
  );
  InMux inmux_21_10_83943_84007 (
    .I(net_83943),
    .O(net_84007)
  );
  CEMux inmux_21_10_83945_84022 (
    .I(net_83945),
    .O(net_84022)
  );
  InMux inmux_21_10_83946_84006 (
    .I(net_83946),
    .O(net_84006)
  );
  InMux inmux_21_10_83947_83978 (
    .I(net_83947),
    .O(net_83978)
  );
  SRMux inmux_21_10_83956_84024 (
    .I(net_83956),
    .O(net_84024)
  );
  InMux inmux_21_10_83963_83976 (
    .I(net_83963),
    .O(net_83976)
  );
  InMux inmux_21_10_83964_83982 (
    .I(net_83964),
    .O(net_83982)
  );
  InMux inmux_21_10_83967_84001 (
    .I(net_83967),
    .O(net_84001)
  );
  InMux inmux_21_10_83972_83985 (
    .I(net_83972),
    .O(net_83985)
  );
  InMux inmux_21_10_83972_84002 (
    .I(net_83972),
    .O(net_84002)
  );
  InMux inmux_21_10_83972_84009 (
    .I(net_83972),
    .O(net_84009)
  );
  ClkMux inmux_21_12_5_84269 (
    .I(net_5),
    .O(net_84269)
  );
  InMux inmux_21_12_84189_84253 (
    .I(net_84189),
    .O(net_84253)
  );
  InMux inmux_21_12_84196_84252 (
    .I(net_84196),
    .O(net_84252)
  );
  InMux inmux_21_12_84197_84254 (
    .I(net_84197),
    .O(net_84254)
  );
  InMux inmux_21_12_84202_84267 (
    .I(net_84202),
    .O(net_84267)
  );
  InMux inmux_21_12_84204_84255 (
    .I(net_84204),
    .O(net_84255)
  );
  InMux inmux_21_12_84217_84235 (
    .I(net_84217),
    .O(net_84235)
  );
  CEMux inmux_21_13_10_84391 (
    .I(net_10),
    .O(net_84391)
  );
  SRMux inmux_21_13_11_84393 (
    .I(net_11),
    .O(net_84393)
  );
  ClkMux inmux_21_13_5_84392 (
    .I(net_5),
    .O(net_84392)
  );
  InMux inmux_21_13_84313_84370 (
    .I(net_84313),
    .O(net_84370)
  );
  InMux inmux_21_13_84314_84381 (
    .I(net_84314),
    .O(net_84381)
  );
  InMux inmux_21_13_84316_84347 (
    .I(net_84316),
    .O(net_84347)
  );
  InMux inmux_21_13_84316_84366 (
    .I(net_84316),
    .O(net_84366)
  );
  InMux inmux_21_13_84316_84371 (
    .I(net_84316),
    .O(net_84371)
  );
  InMux inmux_21_13_84316_84383 (
    .I(net_84316),
    .O(net_84383)
  );
  InMux inmux_21_13_84316_84390 (
    .I(net_84316),
    .O(net_84390)
  );
  InMux inmux_21_13_84319_84353 (
    .I(net_84319),
    .O(net_84353)
  );
  InMux inmux_21_13_84321_84359 (
    .I(net_84321),
    .O(net_84359)
  );
  InMux inmux_21_13_84322_84358 (
    .I(net_84322),
    .O(net_84358)
  );
  InMux inmux_21_13_84324_84351 (
    .I(net_84324),
    .O(net_84351)
  );
  InMux inmux_21_13_84325_84357 (
    .I(net_84325),
    .O(net_84357)
  );
  InMux inmux_21_13_84326_84387 (
    .I(net_84326),
    .O(net_84387)
  );
  InMux inmux_21_13_84327_84369 (
    .I(net_84327),
    .O(net_84369)
  );
  InMux inmux_21_13_84328_84345 (
    .I(net_84328),
    .O(net_84345)
  );
  InMux inmux_21_13_84333_84360 (
    .I(net_84333),
    .O(net_84360)
  );
  InMux inmux_21_13_84334_84352 (
    .I(net_84334),
    .O(net_84352)
  );
  InMux inmux_21_13_84335_84382 (
    .I(net_84335),
    .O(net_84382)
  );
  InMux inmux_21_13_84338_84346 (
    .I(net_84338),
    .O(net_84346)
  );
  InMux inmux_21_13_84341_84364 (
    .I(net_84341),
    .O(net_84364)
  );
  InMux inmux_21_13_84342_84363 (
    .I(net_84342),
    .O(net_84363)
  );
  InMux inmux_21_13_84343_84388 (
    .I(net_84343),
    .O(net_84388)
  );
  ClkMux inmux_21_14_5_84515 (
    .I(net_5),
    .O(net_84515)
  );
  InMux inmux_21_14_84436_84481 (
    .I(net_84436),
    .O(net_84481)
  );
  InMux inmux_21_14_84436_84488 (
    .I(net_84436),
    .O(net_84488)
  );
  InMux inmux_21_14_84437_84489 (
    .I(net_84437),
    .O(net_84489)
  );
  InMux inmux_21_14_84438_84512 (
    .I(net_84438),
    .O(net_84512)
  );
  InMux inmux_21_14_84439_84468 (
    .I(net_84439),
    .O(net_84468)
  );
  InMux inmux_21_14_84439_84477 (
    .I(net_84439),
    .O(net_84477)
  );
  InMux inmux_21_14_84439_84494 (
    .I(net_84439),
    .O(net_84494)
  );
  InMux inmux_21_14_84439_84499 (
    .I(net_84439),
    .O(net_84499)
  );
  InMux inmux_21_14_84439_84504 (
    .I(net_84439),
    .O(net_84504)
  );
  InMux inmux_21_14_84439_84513 (
    .I(net_84439),
    .O(net_84513)
  );
  InMux inmux_21_14_84441_84487 (
    .I(net_84441),
    .O(net_84487)
  );
  InMux inmux_21_14_84442_84505 (
    .I(net_84442),
    .O(net_84505)
  );
  InMux inmux_21_14_84443_84493 (
    .I(net_84443),
    .O(net_84493)
  );
  InMux inmux_21_14_84444_84480 (
    .I(net_84444),
    .O(net_84480)
  );
  InMux inmux_21_14_84445_84500 (
    .I(net_84445),
    .O(net_84500)
  );
  InMux inmux_21_14_84446_84506 (
    .I(net_84446),
    .O(net_84506)
  );
  InMux inmux_21_14_84447_84510 (
    .I(net_84447),
    .O(net_84510)
  );
  InMux inmux_21_14_84448_84475 (
    .I(net_84448),
    .O(net_84475)
  );
  InMux inmux_21_14_84450_84511 (
    .I(net_84450),
    .O(net_84511)
  );
  InMux inmux_21_14_84452_84507 (
    .I(net_84452),
    .O(net_84507)
  );
  InMux inmux_21_14_84453_84501 (
    .I(net_84453),
    .O(net_84501)
  );
  InMux inmux_21_14_84454_84483 (
    .I(net_84454),
    .O(net_84483)
  );
  InMux inmux_21_14_84455_84482 (
    .I(net_84455),
    .O(net_84482)
  );
  InMux inmux_21_14_84456_84476 (
    .I(net_84456),
    .O(net_84476)
  );
  InMux inmux_21_14_84458_84486 (
    .I(net_84458),
    .O(net_84486)
  );
  InMux inmux_21_14_84459_84495 (
    .I(net_84459),
    .O(net_84495)
  );
  CEMux inmux_21_14_84462_84514 (
    .I(net_84462),
    .O(net_84514)
  );
  InMux inmux_21_14_84463_84474 (
    .I(net_84463),
    .O(net_84474)
  );
  InMux inmux_21_14_84465_84498 (
    .I(net_84465),
    .O(net_84498)
  );
  InMux inmux_21_14_84466_84492 (
    .I(net_84466),
    .O(net_84492)
  );
  ClkMux inmux_21_15_5_84638 (
    .I(net_5),
    .O(net_84638)
  );
  InMux inmux_21_15_84558_84610 (
    .I(net_84558),
    .O(net_84610)
  );
  CEMux inmux_21_15_84560_84637 (
    .I(net_84560),
    .O(net_84637)
  );
  InMux inmux_21_15_84561_84609 (
    .I(net_84561),
    .O(net_84609)
  );
  InMux inmux_21_15_84562_84612 (
    .I(net_84562),
    .O(net_84612)
  );
  InMux inmux_21_15_84562_84617 (
    .I(net_84562),
    .O(net_84617)
  );
  InMux inmux_21_15_84562_84629 (
    .I(net_84562),
    .O(net_84629)
  );
  InMux inmux_21_15_84563_84618 (
    .I(net_84563),
    .O(net_84618)
  );
  InMux inmux_21_15_84564_84591 (
    .I(net_84564),
    .O(net_84591)
  );
  InMux inmux_21_15_84566_84621 (
    .I(net_84566),
    .O(net_84621)
  );
  InMux inmux_21_15_84567_84600 (
    .I(net_84567),
    .O(net_84600)
  );
  InMux inmux_21_15_84568_84630 (
    .I(net_84568),
    .O(net_84630)
  );
  InMux inmux_21_15_84569_84593 (
    .I(net_84569),
    .O(net_84593)
  );
  InMux inmux_21_15_84570_84597 (
    .I(net_84570),
    .O(net_84597)
  );
  SRMux inmux_21_15_84571_84639 (
    .I(net_84571),
    .O(net_84639)
  );
  InMux inmux_21_15_84572_84628 (
    .I(net_84572),
    .O(net_84628)
  );
  InMux inmux_21_15_84573_84598 (
    .I(net_84573),
    .O(net_84598)
  );
  InMux inmux_21_15_84573_84603 (
    .I(net_84573),
    .O(net_84603)
  );
  InMux inmux_21_15_84573_84622 (
    .I(net_84573),
    .O(net_84622)
  );
  InMux inmux_21_15_84573_84627 (
    .I(net_84573),
    .O(net_84627)
  );
  InMux inmux_21_15_84573_84636 (
    .I(net_84573),
    .O(net_84636)
  );
  InMux inmux_21_15_84575_84635 (
    .I(net_84575),
    .O(net_84635)
  );
  InMux inmux_21_15_84578_84624 (
    .I(net_84578),
    .O(net_84624)
  );
  InMux inmux_21_15_84581_84604 (
    .I(net_84581),
    .O(net_84604)
  );
  InMux inmux_21_15_84582_84592 (
    .I(net_84582),
    .O(net_84592)
  );
  InMux inmux_21_15_84582_84599 (
    .I(net_84582),
    .O(net_84599)
  );
  InMux inmux_21_15_84582_84633 (
    .I(net_84582),
    .O(net_84633)
  );
  InMux inmux_21_15_84583_84615 (
    .I(net_84583),
    .O(net_84615)
  );
  InMux inmux_21_15_84584_84594 (
    .I(net_84584),
    .O(net_84594)
  );
  InMux inmux_21_15_84585_84605 (
    .I(net_84585),
    .O(net_84605)
  );
  InMux inmux_21_15_84586_84623 (
    .I(net_84586),
    .O(net_84623)
  );
  InMux inmux_21_15_84589_84634 (
    .I(net_84589),
    .O(net_84634)
  );
  CEMux inmux_21_16_10_84760 (
    .I(net_10),
    .O(net_84760)
  );
  ClkMux inmux_21_16_5_84761 (
    .I(net_5),
    .O(net_84761)
  );
  InMux inmux_21_16_84682_84732 (
    .I(net_84682),
    .O(net_84732)
  );
  InMux inmux_21_16_84686_84739 (
    .I(net_84686),
    .O(net_84739)
  );
  InMux inmux_21_16_84694_84750 (
    .I(net_84694),
    .O(net_84750)
  );
  InMux inmux_21_16_84696_84735 (
    .I(net_84696),
    .O(net_84735)
  );
  InMux inmux_21_16_84698_84741 (
    .I(net_84698),
    .O(net_84741)
  );
  InMux inmux_21_16_84706_84733 (
    .I(net_84706),
    .O(net_84733)
  );
  InMux inmux_21_16_84711_84734 (
    .I(net_84711),
    .O(net_84734)
  );
  ClkMux inmux_21_17_5_84884 (
    .I(net_5),
    .O(net_84884)
  );
  InMux inmux_21_17_84806_84875 (
    .I(net_84806),
    .O(net_84875)
  );
  InMux inmux_21_17_84808_84870 (
    .I(net_84808),
    .O(net_84870)
  );
  InMux inmux_21_17_84812_84876 (
    .I(net_84812),
    .O(net_84876)
  );
  InMux inmux_21_17_84813_84873 (
    .I(net_84813),
    .O(net_84873)
  );
  InMux inmux_21_17_84814_84874 (
    .I(net_84814),
    .O(net_84874)
  );
  InMux inmux_21_17_84815_84837 (
    .I(net_84815),
    .O(net_84837)
  );
  InMux inmux_21_17_84817_84839 (
    .I(net_84817),
    .O(net_84839)
  );
  InMux inmux_21_17_84821_84850 (
    .I(net_84821),
    .O(net_84850)
  );
  InMux inmux_21_17_84822_84882 (
    .I(net_84822),
    .O(net_84882)
  );
  InMux inmux_21_17_84824_84846 (
    .I(net_84824),
    .O(net_84846)
  );
  InMux inmux_21_17_84825_84845 (
    .I(net_84825),
    .O(net_84845)
  );
  InMux inmux_21_17_84826_84858 (
    .I(net_84826),
    .O(net_84858)
  );
  InMux inmux_21_17_84827_84843 (
    .I(net_84827),
    .O(net_84843)
  );
  InMux inmux_21_17_84829_84851 (
    .I(net_84829),
    .O(net_84851)
  );
  InMux inmux_21_17_84830_84852 (
    .I(net_84830),
    .O(net_84852)
  );
  InMux inmux_21_17_84831_84844 (
    .I(net_84831),
    .O(net_84844)
  );
  InMux inmux_21_17_84832_84838 (
    .I(net_84832),
    .O(net_84838)
  );
  InMux inmux_21_17_84833_84863 (
    .I(net_84833),
    .O(net_84863)
  );
  InMux inmux_21_17_84834_84840 (
    .I(net_84834),
    .O(net_84840)
  );
  InMux inmux_21_17_84835_84849 (
    .I(net_84835),
    .O(net_84849)
  );
  CEMux inmux_21_18_10_85006 (
    .I(net_10),
    .O(net_85006)
  );
  ClkMux inmux_21_18_5_85007 (
    .I(net_5),
    .O(net_85007)
  );
  InMux inmux_21_18_84928_84985 (
    .I(net_84928),
    .O(net_84985)
  );
  InMux inmux_21_18_84929_84984 (
    .I(net_84929),
    .O(net_84984)
  );
  InMux inmux_21_18_84930_84975 (
    .I(net_84930),
    .O(net_84975)
  );
  InMux inmux_21_18_84931_84972 (
    .I(net_84931),
    .O(net_84972)
  );
  InMux inmux_21_18_84935_84992 (
    .I(net_84935),
    .O(net_84992)
  );
  InMux inmux_21_18_84935_85002 (
    .I(net_84935),
    .O(net_85002)
  );
  InMux inmux_21_18_84936_84996 (
    .I(net_84936),
    .O(net_84996)
  );
  InMux inmux_21_18_84938_85003 (
    .I(net_84938),
    .O(net_85003)
  );
  InMux inmux_21_18_84939_84997 (
    .I(net_84939),
    .O(net_84997)
  );
  InMux inmux_21_18_84940_84991 (
    .I(net_84940),
    .O(net_84991)
  );
  InMux inmux_21_18_84940_85005 (
    .I(net_84940),
    .O(net_85005)
  );
  InMux inmux_21_18_84941_84963 (
    .I(net_84941),
    .O(net_84963)
  );
  InMux inmux_21_18_84941_84966 (
    .I(net_84941),
    .O(net_84966)
  );
  InMux inmux_21_18_84941_84980 (
    .I(net_84941),
    .O(net_84980)
  );
  InMux inmux_21_18_84952_84993 (
    .I(net_84952),
    .O(net_84993)
  );
  InMux inmux_21_18_84953_84973 (
    .I(net_84953),
    .O(net_84973)
  );
  InMux inmux_21_18_84953_84987 (
    .I(net_84953),
    .O(net_84987)
  );
  InMux inmux_21_18_84953_84999 (
    .I(net_84953),
    .O(net_84999)
  );
  InMux inmux_21_18_84955_85004 (
    .I(net_84955),
    .O(net_85004)
  );
  InMux inmux_21_18_84957_84990 (
    .I(net_84957),
    .O(net_84990)
  );
  CEMux inmux_21_19_10_85129 (
    .I(net_10),
    .O(net_85129)
  );
  ClkMux inmux_21_19_5_85130 (
    .I(net_5),
    .O(net_85130)
  );
  InMux inmux_21_19_85064_85098 (
    .I(net_85064),
    .O(net_85098)
  );
  InMux inmux_21_19_85064_85103 (
    .I(net_85064),
    .O(net_85103)
  );
  InMux inmux_21_6_83456_83504 (
    .I(net_83456),
    .O(net_83504)
  );
  InMux inmux_21_6_83456_83514 (
    .I(net_83456),
    .O(net_83514)
  );
  InMux inmux_21_6_83460_83503 (
    .I(net_83460),
    .O(net_83503)
  );
  InMux inmux_21_6_83466_83505 (
    .I(net_83466),
    .O(net_83505)
  );
  InMux inmux_21_6_83466_83515 (
    .I(net_83466),
    .O(net_83515)
  );
  ClkMux inmux_21_9_5_83900 (
    .I(net_5),
    .O(net_83900)
  );
  CEMux inmux_21_9_83822_83899 (
    .I(net_83822),
    .O(net_83899)
  );
  InMux inmux_21_9_83828_83854 (
    .I(net_83828),
    .O(net_83854)
  );
  InMux inmux_21_9_83828_83892 (
    .I(net_83828),
    .O(net_83892)
  );
  InMux inmux_21_9_83833_83867 (
    .I(net_83833),
    .O(net_83867)
  );
  InMux inmux_21_9_83833_83889 (
    .I(net_83833),
    .O(net_83889)
  );
  InMux inmux_21_9_83835_83855 (
    .I(net_83835),
    .O(net_83855)
  );
  InMux inmux_21_9_83843_83866 (
    .I(net_83843),
    .O(net_83866)
  );
  InMux inmux_21_9_83843_83890 (
    .I(net_83843),
    .O(net_83890)
  );
  SRMux inmux_21_9_83849_83901 (
    .I(net_83849),
    .O(net_83901)
  );
  IoInMux inmux_22_0_86579_86563 (
    .I(net_86579),
    .O(net_86563)
  );
  ClkMux inmux_22_13_5_88223 (
    .I(net_5),
    .O(net_88223)
  );
  InMux inmux_22_13_88152_88190 (
    .I(net_88152),
    .O(net_88190)
  );
  InMux inmux_22_13_88166_88208 (
    .I(net_88166),
    .O(net_88208)
  );
  CEMux inmux_22_14_10_88345 (
    .I(net_10),
    .O(net_88345)
  );
  SRMux inmux_22_14_11_88347 (
    .I(net_11),
    .O(net_88347)
  );
  ClkMux inmux_22_14_5_88346 (
    .I(net_5),
    .O(net_88346)
  );
  InMux inmux_22_14_88270_88318 (
    .I(net_88270),
    .O(net_88318)
  );
  InMux inmux_22_14_88278_88319 (
    .I(net_88278),
    .O(net_88319)
  );
  InMux inmux_22_14_88279_88320 (
    .I(net_88279),
    .O(net_88320)
  );
  ClkMux inmux_22_15_5_88469 (
    .I(net_5),
    .O(net_88469)
  );
  InMux inmux_22_15_88417_88449 (
    .I(net_88417),
    .O(net_88449)
  );
  InMux inmux_22_15_88419_88437 (
    .I(net_88419),
    .O(net_88437)
  );
  CEMux inmux_22_16_10_88591 (
    .I(net_10),
    .O(net_88591)
  );
  SRMux inmux_22_16_11_88593 (
    .I(net_11),
    .O(net_88593)
  );
  ClkMux inmux_22_16_5_88592 (
    .I(net_5),
    .O(net_88592)
  );
  InMux inmux_22_16_88534_88588 (
    .I(net_88534),
    .O(net_88588)
  );
  InMux inmux_22_16_88539_88590 (
    .I(net_88539),
    .O(net_88590)
  );
  InMux inmux_22_17_88636_88693 (
    .I(net_88636),
    .O(net_88693)
  );
  InMux inmux_22_17_88638_88705 (
    .I(net_88638),
    .O(net_88705)
  );
  InMux inmux_22_17_88639_88699 (
    .I(net_88639),
    .O(net_88699)
  );
  InMux inmux_22_17_88640_88669 (
    .I(net_88640),
    .O(net_88669)
  );
  InMux inmux_22_17_88642_88681 (
    .I(net_88642),
    .O(net_88681)
  );
  InMux inmux_22_17_88646_88687 (
    .I(net_88646),
    .O(net_88687)
  );
  InMux inmux_22_17_88647_88676 (
    .I(net_88647),
    .O(net_88676)
  );
  InMux inmux_22_17_88650_88670 (
    .I(net_88650),
    .O(net_88670)
  );
  InMux inmux_22_17_88656_88712 (
    .I(net_88656),
    .O(net_88712)
  );
  InMux inmux_22_17_88667_88677 (
    .I(net_88667),
    .O(net_88677)
  );
  InMux inmux_22_17_88673_88683 (
    .I(net_88673),
    .O(net_88683)
  );
  InMux inmux_22_17_88679_88689 (
    .I(net_88679),
    .O(net_88689)
  );
  InMux inmux_22_17_88685_88695 (
    .I(net_88685),
    .O(net_88695)
  );
  InMux inmux_22_17_88691_88701 (
    .I(net_88691),
    .O(net_88701)
  );
  InMux inmux_22_17_88697_88707 (
    .I(net_88697),
    .O(net_88707)
  );
  InMux inmux_22_17_88703_88713 (
    .I(net_88703),
    .O(net_88713)
  );
  ClkMux inmux_22_9_5_87731 (
    .I(net_5),
    .O(net_87731)
  );
  InMux inmux_22_9_87652_87692 (
    .I(net_87652),
    .O(net_87692)
  );
  SRMux inmux_22_9_87655_87732 (
    .I(net_87655),
    .O(net_87732)
  );
  CEMux inmux_22_9_87669_87730 (
    .I(net_87669),
    .O(net_87730)
  );
  ClkMux inmux_23_9_5_91562 (
    .I(net_5),
    .O(net_91562)
  );
  InMux inmux_23_9_91484_91529 (
    .I(net_91484),
    .O(net_91529)
  );
  InMux inmux_23_9_91484_91558 (
    .I(net_91484),
    .O(net_91558)
  );
  InMux inmux_23_9_91491_91522 (
    .I(net_91491),
    .O(net_91522)
  );
  InMux inmux_23_9_91491_91560 (
    .I(net_91491),
    .O(net_91560)
  );
  CEMux inmux_23_9_91493_91561 (
    .I(net_91493),
    .O(net_91561)
  );
  SRMux inmux_23_9_91495_91563 (
    .I(net_91495),
    .O(net_91563)
  );
  InMux inmux_23_9_91506_91516 (
    .I(net_91506),
    .O(net_91516)
  );
  InMux inmux_23_9_91506_91557 (
    .I(net_91506),
    .O(net_91557)
  );
  InMux inmux_23_9_91520_91530 (
    .I(net_91520),
    .O(net_91530)
  );
  InMux inmux_2_19_13545_13558 (
    .I(net_13545),
    .O(net_13558)
  );
  InMux inmux_2_19_13551_13561 (
    .I(net_13551),
    .O(net_13561)
  );
  InMux inmux_2_19_13554_13560 (
    .I(net_13554),
    .O(net_13560)
  );
  InMux inmux_2_19_13555_13559 (
    .I(net_13555),
    .O(net_13559)
  );
  InMux inmux_2_8_12178_12248 (
    .I(net_12178),
    .O(net_12248)
  );
  InMux inmux_2_8_12179_12206 (
    .I(net_12179),
    .O(net_12206)
  );
  InMux inmux_2_8_12179_12247 (
    .I(net_12179),
    .O(net_12247)
  );
  SRMux inmux_2_8_12185_12253 (
    .I(net_12185),
    .O(net_12253)
  );
  InMux inmux_2_8_12191_12225 (
    .I(net_12191),
    .O(net_12225)
  );
  InMux inmux_2_8_12191_12249 (
    .I(net_12191),
    .O(net_12249)
  );
  InMux inmux_2_8_12192_12231 (
    .I(net_12192),
    .O(net_12231)
  );
  InMux inmux_2_8_12192_12241 (
    .I(net_12192),
    .O(net_12241)
  );
  InMux inmux_2_8_12198_12218 (
    .I(net_12198),
    .O(net_12218)
  );
  InMux inmux_2_8_12198_12244 (
    .I(net_12198),
    .O(net_12244)
  );
  InMux inmux_2_8_12200_12213 (
    .I(net_12200),
    .O(net_12213)
  );
  InMux inmux_2_8_12200_12242 (
    .I(net_12200),
    .O(net_12242)
  );
  InMux inmux_2_8_12201_12236 (
    .I(net_12201),
    .O(net_12236)
  );
  InMux inmux_2_8_12201_12243 (
    .I(net_12201),
    .O(net_12243)
  );
  InMux inmux_2_8_12210_12220 (
    .I(net_12210),
    .O(net_12220)
  );
  InMux inmux_2_8_12216_12226 (
    .I(net_12216),
    .O(net_12226)
  );
  InMux inmux_2_8_12222_12232 (
    .I(net_12222),
    .O(net_12232)
  );
  InMux inmux_2_8_12228_12238 (
    .I(net_12228),
    .O(net_12238)
  );
  ClkMux inmux_2_8_5_12252 (
    .I(net_5),
    .O(net_12252)
  );
  InMux inmux_3_13_16620_16665 (
    .I(net_16620),
    .O(net_16665)
  );
  InMux inmux_3_13_16620_16689 (
    .I(net_16620),
    .O(net_16689)
  );
  InMux inmux_3_13_16628_16659 (
    .I(net_16628),
    .O(net_16659)
  );
  InMux inmux_3_13_16628_16688 (
    .I(net_16628),
    .O(net_16688)
  );
  SRMux inmux_3_13_16631_16699 (
    .I(net_16631),
    .O(net_16699)
  );
  InMux inmux_3_13_16632_16695 (
    .I(net_16632),
    .O(net_16695)
  );
  InMux inmux_3_13_16639_16652 (
    .I(net_16639),
    .O(net_16652)
  );
  InMux inmux_3_13_16639_16693 (
    .I(net_16639),
    .O(net_16693)
  );
  InMux inmux_3_13_16645_16670 (
    .I(net_16645),
    .O(net_16670)
  );
  InMux inmux_3_13_16645_16694 (
    .I(net_16645),
    .O(net_16694)
  );
  InMux inmux_3_13_16646_16676 (
    .I(net_16646),
    .O(net_16676)
  );
  InMux inmux_3_13_16646_16690 (
    .I(net_16646),
    .O(net_16690)
  );
  InMux inmux_3_13_16647_16682 (
    .I(net_16647),
    .O(net_16682)
  );
  InMux inmux_3_13_16647_16687 (
    .I(net_16647),
    .O(net_16687)
  );
  InMux inmux_3_13_16656_16666 (
    .I(net_16656),
    .O(net_16666)
  );
  InMux inmux_3_13_16662_16672 (
    .I(net_16662),
    .O(net_16672)
  );
  InMux inmux_3_13_16668_16678 (
    .I(net_16668),
    .O(net_16678)
  );
  InMux inmux_3_13_16674_16684 (
    .I(net_16674),
    .O(net_16684)
  );
  ClkMux inmux_3_13_5_16698 (
    .I(net_5),
    .O(net_16698)
  );
  InMux inmux_3_14_16759_16786 (
    .I(net_16759),
    .O(net_16786)
  );
  CEMux inmux_3_14_16768_16820 (
    .I(net_16768),
    .O(net_16820)
  );
  SRMux inmux_3_14_16770_16822 (
    .I(net_16770),
    .O(net_16822)
  );
  ClkMux inmux_3_14_5_16821 (
    .I(net_5),
    .O(net_16821)
  );
  InMux inmux_3_18_17237_17292 (
    .I(net_17237),
    .O(net_17292)
  );
  InMux inmux_3_18_17238_17298 (
    .I(net_17238),
    .O(net_17298)
  );
  InMux inmux_3_18_17239_17304 (
    .I(net_17239),
    .O(net_17304)
  );
  InMux inmux_3_18_17242_17273 (
    .I(net_17242),
    .O(net_17273)
  );
  InMux inmux_3_18_17251_17280 (
    .I(net_17251),
    .O(net_17280)
  );
  InMux inmux_3_18_17252_17286 (
    .I(net_17252),
    .O(net_17286)
  );
  InMux inmux_3_18_17256_17267 (
    .I(net_17256),
    .O(net_17267)
  );
  InMux inmux_3_18_17264_17309 (
    .I(net_17264),
    .O(net_17309)
  );
  InMux inmux_3_18_17271_17281 (
    .I(net_17271),
    .O(net_17281)
  );
  InMux inmux_3_18_17277_17287 (
    .I(net_17277),
    .O(net_17287)
  );
  InMux inmux_3_18_17283_17293 (
    .I(net_17283),
    .O(net_17293)
  );
  InMux inmux_3_18_17289_17299 (
    .I(net_17289),
    .O(net_17299)
  );
  InMux inmux_3_18_17295_17305 (
    .I(net_17295),
    .O(net_17305)
  );
  InMux inmux_3_18_17301_17311 (
    .I(net_17301),
    .O(net_17311)
  );
  ClkMux inmux_3_18_5_17313 (
    .I(net_5),
    .O(net_17313)
  );
  InMux inmux_3_19_17351_17392 (
    .I(net_17351),
    .O(net_17392)
  );
  InMux inmux_3_19_17357_17397 (
    .I(net_17357),
    .O(net_17397)
  );
  InMux inmux_3_19_17362_17427 (
    .I(net_17362),
    .O(net_17427)
  );
  InMux inmux_3_19_17364_17390 (
    .I(net_17364),
    .O(net_17390)
  );
  InMux inmux_3_19_17367_17408 (
    .I(net_17367),
    .O(net_17408)
  );
  InMux inmux_3_19_17376_17415 (
    .I(net_17376),
    .O(net_17415)
  );
  InMux inmux_3_19_17377_17421 (
    .I(net_17377),
    .O(net_17421)
  );
  InMux inmux_3_19_17379_17433 (
    .I(net_17379),
    .O(net_17433)
  );
  InMux inmux_3_19_17382_17402 (
    .I(net_17382),
    .O(net_17402)
  );
  InMux inmux_3_19_17388_17398 (
    .I(net_17388),
    .O(net_17398)
  );
  InMux inmux_3_19_17394_17404 (
    .I(net_17394),
    .O(net_17404)
  );
  InMux inmux_3_19_17400_17410 (
    .I(net_17400),
    .O(net_17410)
  );
  InMux inmux_3_19_17406_17416 (
    .I(net_17406),
    .O(net_17416)
  );
  InMux inmux_3_19_17412_17422 (
    .I(net_17412),
    .O(net_17422)
  );
  InMux inmux_3_19_17418_17428 (
    .I(net_17418),
    .O(net_17428)
  );
  InMux inmux_3_19_17424_17434 (
    .I(net_17424),
    .O(net_17434)
  );
  ClkMux inmux_3_19_5_17436 (
    .I(net_5),
    .O(net_17436)
  );
  InMux inmux_3_20_17474_17515 (
    .I(net_17474),
    .O(net_17515)
  );
  InMux inmux_3_20_17481_17526 (
    .I(net_17481),
    .O(net_17526)
  );
  InMux inmux_3_20_17493_17549 (
    .I(net_17493),
    .O(net_17549)
  );
  InMux inmux_3_20_17495_17514 (
    .I(net_17495),
    .O(net_17514)
  );
  InMux inmux_3_20_17500_17544 (
    .I(net_17500),
    .O(net_17544)
  );
  InMux inmux_3_20_17504_17519 (
    .I(net_17504),
    .O(net_17519)
  );
  InMux inmux_3_20_17506_17531 (
    .I(net_17506),
    .O(net_17531)
  );
  InMux inmux_3_20_17507_17537 (
    .I(net_17507),
    .O(net_17537)
  );
  InMux inmux_3_20_17510_17555 (
    .I(net_17510),
    .O(net_17555)
  );
  InMux inmux_3_20_17511_17521 (
    .I(net_17511),
    .O(net_17521)
  );
  InMux inmux_3_20_17517_17527 (
    .I(net_17517),
    .O(net_17527)
  );
  InMux inmux_3_20_17523_17533 (
    .I(net_17523),
    .O(net_17533)
  );
  InMux inmux_3_20_17529_17539 (
    .I(net_17529),
    .O(net_17539)
  );
  InMux inmux_3_20_17535_17545 (
    .I(net_17535),
    .O(net_17545)
  );
  InMux inmux_3_20_17541_17551 (
    .I(net_17541),
    .O(net_17551)
  );
  InMux inmux_3_20_17547_17557 (
    .I(net_17547),
    .O(net_17557)
  );
  ClkMux inmux_3_20_5_17559 (
    .I(net_5),
    .O(net_17559)
  );
  InMux inmux_3_7_15887_15955 (
    .I(net_15887),
    .O(net_15955)
  );
  SRMux inmux_3_7_15893_15961 (
    .I(net_15893),
    .O(net_15961)
  );
  InMux inmux_3_7_15895_15958 (
    .I(net_15895),
    .O(net_15958)
  );
  ClkMux inmux_3_7_5_15960 (
    .I(net_5),
    .O(net_15960)
  );
  CEMux inmux_3_8_16014_16082 (
    .I(net_16014),
    .O(net_16082)
  );
  InMux inmux_3_8_16015_16061 (
    .I(net_16015),
    .O(net_16061)
  );
  SRMux inmux_3_8_16016_16084 (
    .I(net_16016),
    .O(net_16084)
  );
  ClkMux inmux_3_8_5_16083 (
    .I(net_5),
    .O(net_16083)
  );
  InMux inmux_4_12_20341_20371 (
    .I(net_20341),
    .O(net_20371)
  );
  InMux inmux_4_12_20352_20374 (
    .I(net_20352),
    .O(net_20374)
  );
  ClkMux inmux_4_12_5_20406 (
    .I(net_5),
    .O(net_20406)
  );
  InMux inmux_4_13_20461_20514 (
    .I(net_20461),
    .O(net_20514)
  );
  SRMux inmux_4_13_20462_20530 (
    .I(net_20462),
    .O(net_20530)
  );
  InMux inmux_4_13_20478_20513 (
    .I(net_20478),
    .O(net_20513)
  );
  ClkMux inmux_4_13_5_20529 (
    .I(net_5),
    .O(net_20529)
  );
  InMux inmux_4_17_20942_20982 (
    .I(net_20942),
    .O(net_20982)
  );
  CEMux inmux_4_17_20968_21020 (
    .I(net_20968),
    .O(net_21020)
  );
  ClkMux inmux_4_17_5_21021 (
    .I(net_5),
    .O(net_21021)
  );
  InMux inmux_4_18_21065_21098 (
    .I(net_21065),
    .O(net_21098)
  );
  InMux inmux_4_18_21066_21097 (
    .I(net_21066),
    .O(net_21097)
  );
  InMux inmux_4_18_21069_21136 (
    .I(net_21069),
    .O(net_21136)
  );
  InMux inmux_4_18_21070_21135 (
    .I(net_21070),
    .O(net_21135)
  );
  InMux inmux_4_18_21072_21112 (
    .I(net_21072),
    .O(net_21112)
  );
  InMux inmux_4_18_21073_21109 (
    .I(net_21073),
    .O(net_21109)
  );
  InMux inmux_4_18_21075_21099 (
    .I(net_21075),
    .O(net_21099)
  );
  InMux inmux_4_18_21076_21134 (
    .I(net_21076),
    .O(net_21134)
  );
  InMux inmux_4_18_21078_21141 (
    .I(net_21078),
    .O(net_21141)
  );
  InMux inmux_4_18_21086_21111 (
    .I(net_21086),
    .O(net_21111)
  );
  InMux inmux_4_18_21087_21100 (
    .I(net_21087),
    .O(net_21100)
  );
  InMux inmux_4_18_21087_21139 (
    .I(net_21087),
    .O(net_21139)
  );
  InMux inmux_4_18_21089_21133 (
    .I(net_21089),
    .O(net_21133)
  );
  ClkMux inmux_4_18_5_21144 (
    .I(net_5),
    .O(net_21144)
  );
  InMux inmux_4_19_21189_21229 (
    .I(net_21189),
    .O(net_21229)
  );
  InMux inmux_4_19_21190_21233 (
    .I(net_21190),
    .O(net_21233)
  );
  InMux inmux_4_19_21195_21247 (
    .I(net_21195),
    .O(net_21247)
  );
  InMux inmux_4_19_21196_21227 (
    .I(net_21196),
    .O(net_21227)
  );
  InMux inmux_4_19_21197_21235 (
    .I(net_21197),
    .O(net_21235)
  );
  InMux inmux_4_19_21199_21228 (
    .I(net_21199),
    .O(net_21228)
  );
  InMux inmux_4_19_21202_21232 (
    .I(net_21202),
    .O(net_21232)
  );
  InMux inmux_4_19_21203_21234 (
    .I(net_21203),
    .O(net_21234)
  );
  InMux inmux_4_19_21210_21245 (
    .I(net_21210),
    .O(net_21245)
  );
  InMux inmux_4_19_21211_21226 (
    .I(net_21211),
    .O(net_21226)
  );
  InMux inmux_4_19_21216_21246 (
    .I(net_21216),
    .O(net_21246)
  );
  InMux inmux_4_19_21218_21244 (
    .I(net_21218),
    .O(net_21244)
  );
  InMux inmux_4_20_21313_21349 (
    .I(net_21313),
    .O(net_21349)
  );
  InMux inmux_4_20_21316_21352 (
    .I(net_21316),
    .O(net_21352)
  );
  InMux inmux_4_20_21319_21350 (
    .I(net_21319),
    .O(net_21350)
  );
  InMux inmux_4_20_21322_21351 (
    .I(net_21322),
    .O(net_21351)
  );
  CEMux inmux_5_12_24159_24236 (
    .I(net_24159),
    .O(net_24236)
  );
  InMux inmux_5_12_24175_24202 (
    .I(net_24175),
    .O(net_24202)
  );
  ClkMux inmux_5_12_5_24237 (
    .I(net_5),
    .O(net_24237)
  );
  InMux inmux_5_20_25152_25188 (
    .I(net_25152),
    .O(net_25188)
  );
  ClkMux inmux_5_20_5_25221 (
    .I(net_5),
    .O(net_25221)
  );
  CEMux inmux_5_20_8_25220 (
    .I(net_8),
    .O(net_25220)
  );
  InMux inmux_5_5_23327_23331 (
    .I(net_23327),
    .O(net_23331)
  );
  ClkMux inmux_5_5_5_23376 (
    .I(net_5),
    .O(net_23376)
  );
  IoInMux inmux_6_0_26539_26528 (
    .I(net_26539),
    .O(net_26528)
  );
  CEMux inmux_6_0_26547_26534 (
    .I(net_26547),
    .O(net_26534)
  );
  ClkMux inmux_6_0_5_26535 (
    .I(net_5),
    .O(net_26535)
  );
  ClkMux inmux_6_0_5_26536 (
    .I(net_5),
    .O(net_26536)
  );
  IoInMux inmux_7_0_29743_29728 (
    .I(net_29743),
    .O(net_29728)
  );
  CEMux inmux_7_0_29747_29734 (
    .I(net_29747),
    .O(net_29734)
  );
  ClkMux inmux_7_0_5_29735 (
    .I(net_5),
    .O(net_29735)
  );
  ClkMux inmux_7_0_5_29736 (
    .I(net_5),
    .O(net_29736)
  );
  InMux inmux_7_12_31207_31239 (
    .I(net_31207),
    .O(net_31239)
  );
  InMux inmux_7_12_31207_31251 (
    .I(net_31207),
    .O(net_31251)
  );
  InMux inmux_7_12_31208_31228 (
    .I(net_31208),
    .O(net_31228)
  );
  InMux inmux_7_12_31208_31252 (
    .I(net_31208),
    .O(net_31252)
  );
  InMux inmux_7_12_31213_31223 (
    .I(net_31213),
    .O(net_31223)
  );
  InMux inmux_7_12_31213_31254 (
    .I(net_31213),
    .O(net_31254)
  );
  InMux inmux_7_12_31214_31234 (
    .I(net_31214),
    .O(net_31234)
  );
  InMux inmux_7_12_31214_31253 (
    .I(net_31214),
    .O(net_31253)
  );
  InMux inmux_7_12_31226_31236 (
    .I(net_31226),
    .O(net_31236)
  );
  InMux inmux_7_12_31232_31242 (
    .I(net_31232),
    .O(net_31242)
  );
  ClkMux inmux_7_12_5_31268 (
    .I(net_5),
    .O(net_31268)
  );
  InMux inmux_7_1_29814_29836 (
    .I(net_29814),
    .O(net_29836)
  );
  InMux inmux_7_1_29826_29837 (
    .I(net_29826),
    .O(net_29837)
  );
  InMux inmux_8_10_34775_34820 (
    .I(net_34775),
    .O(net_34820)
  );
  InMux inmux_8_10_34775_34842 (
    .I(net_34775),
    .O(net_34842)
  );
  SRMux inmux_8_10_34777_34854 (
    .I(net_34777),
    .O(net_34854)
  );
  InMux inmux_8_10_34778_34838 (
    .I(net_34778),
    .O(net_34838)
  );
  InMux inmux_8_10_34778_34843 (
    .I(net_34778),
    .O(net_34843)
  );
  InMux inmux_8_10_34779_34849 (
    .I(net_34779),
    .O(net_34849)
  );
  InMux inmux_8_10_34786_34813 (
    .I(net_34786),
    .O(net_34813)
  );
  InMux inmux_8_10_34786_34844 (
    .I(net_34786),
    .O(net_34844)
  );
  InMux inmux_8_10_34799_34807 (
    .I(net_34799),
    .O(net_34807)
  );
  InMux inmux_8_10_34799_34850 (
    .I(net_34799),
    .O(net_34850)
  );
  InMux inmux_8_10_34800_34825 (
    .I(net_34800),
    .O(net_34825)
  );
  InMux inmux_8_10_34800_34851 (
    .I(net_34800),
    .O(net_34851)
  );
  InMux inmux_8_10_34801_34831 (
    .I(net_34801),
    .O(net_34831)
  );
  InMux inmux_8_10_34801_34845 (
    .I(net_34801),
    .O(net_34845)
  );
  InMux inmux_8_10_34811_34821 (
    .I(net_34811),
    .O(net_34821)
  );
  InMux inmux_8_10_34817_34827 (
    .I(net_34817),
    .O(net_34827)
  );
  InMux inmux_8_10_34823_34833 (
    .I(net_34823),
    .O(net_34833)
  );
  InMux inmux_8_10_34829_34839 (
    .I(net_34829),
    .O(net_34839)
  );
  ClkMux inmux_8_10_5_34853 (
    .I(net_5),
    .O(net_34853)
  );
  CEMux inmux_8_11_34898_34975 (
    .I(net_34898),
    .O(net_34975)
  );
  InMux inmux_8_11_34901_34961 (
    .I(net_34901),
    .O(net_34961)
  );
  SRMux inmux_8_11_34925_34977 (
    .I(net_34925),
    .O(net_34977)
  );
  ClkMux inmux_8_11_5_34976 (
    .I(net_5),
    .O(net_34976)
  );
  InMux inmux_8_12_35020_35058 (
    .I(net_35020),
    .O(net_35058)
  );
  SRMux inmux_8_12_35023_35100 (
    .I(net_35023),
    .O(net_35100)
  );
  InMux inmux_8_12_35045_35060 (
    .I(net_35045),
    .O(net_35060)
  );
  ClkMux inmux_8_12_5_35099 (
    .I(net_5),
    .O(net_35099)
  );
  InMux inmux_8_17_35651_35699 (
    .I(net_35651),
    .O(net_35699)
  );
  ClkMux inmux_8_17_5_35714 (
    .I(net_5),
    .O(net_35714)
  );
  SRMux inmux_8_23_36376_36453 (
    .I(net_36376),
    .O(net_36453)
  );
  InMux inmux_8_23_36393_36435 (
    .I(net_36393),
    .O(net_36435)
  );
  InMux inmux_8_23_36401_36436 (
    .I(net_36401),
    .O(net_36436)
  );
  ClkMux inmux_8_23_5_36452 (
    .I(net_5),
    .O(net_36452)
  );
  CEMux inmux_8_24_36497_36574 (
    .I(net_36497),
    .O(net_36574)
  );
  SRMux inmux_8_24_36508_36576 (
    .I(net_36508),
    .O(net_36576)
  );
  InMux inmux_8_24_36517_36564 (
    .I(net_36517),
    .O(net_36564)
  );
  ClkMux inmux_8_24_5_36575 (
    .I(net_5),
    .O(net_36575)
  );
  InMux inmux_8_25_36621_36671 (
    .I(net_36621),
    .O(net_36671)
  );
  InMux inmux_8_25_36621_36688 (
    .I(net_36621),
    .O(net_36688)
  );
  SRMux inmux_8_25_36622_36699 (
    .I(net_36622),
    .O(net_36699)
  );
  InMux inmux_8_25_36624_36658 (
    .I(net_36624),
    .O(net_36658)
  );
  InMux inmux_8_25_36624_36696 (
    .I(net_36624),
    .O(net_36696)
  );
  InMux inmux_8_25_36628_36652 (
    .I(net_36628),
    .O(net_36652)
  );
  InMux inmux_8_25_36628_36695 (
    .I(net_36628),
    .O(net_36695)
  );
  InMux inmux_8_25_36630_36676 (
    .I(net_36630),
    .O(net_36676)
  );
  InMux inmux_8_25_36630_36693 (
    .I(net_36630),
    .O(net_36693)
  );
  InMux inmux_8_25_36633_36689 (
    .I(net_36633),
    .O(net_36689)
  );
  InMux inmux_8_25_36636_36665 (
    .I(net_36636),
    .O(net_36665)
  );
  InMux inmux_8_25_36636_36694 (
    .I(net_36636),
    .O(net_36694)
  );
  InMux inmux_8_25_36647_36682 (
    .I(net_36647),
    .O(net_36682)
  );
  InMux inmux_8_25_36647_36687 (
    .I(net_36647),
    .O(net_36687)
  );
  InMux inmux_8_25_36656_36666 (
    .I(net_36656),
    .O(net_36666)
  );
  InMux inmux_8_25_36662_36672 (
    .I(net_36662),
    .O(net_36672)
  );
  InMux inmux_8_25_36668_36678 (
    .I(net_36668),
    .O(net_36678)
  );
  InMux inmux_8_25_36674_36684 (
    .I(net_36674),
    .O(net_36684)
  );
  ClkMux inmux_8_25_5_36698 (
    .I(net_5),
    .O(net_36698)
  );
  InMux inmux_8_2_33791_33831 (
    .I(net_33791),
    .O(net_33831)
  );
  InMux inmux_8_2_33797_33828 (
    .I(net_33797),
    .O(net_33828)
  );
  InMux inmux_8_2_33797_33835 (
    .I(net_33797),
    .O(net_33835)
  );
  InMux inmux_8_2_33802_33843 (
    .I(net_33802),
    .O(net_33843)
  );
  InMux inmux_8_2_33802_33853 (
    .I(net_33802),
    .O(net_33853)
  );
  InMux inmux_8_2_33802_33860 (
    .I(net_33802),
    .O(net_33860)
  );
  InMux inmux_8_2_33802_33865 (
    .I(net_33802),
    .O(net_33865)
  );
  InMux inmux_8_2_33803_33849 (
    .I(net_33803),
    .O(net_33849)
  );
  InMux inmux_8_2_33805_33848 (
    .I(net_33805),
    .O(net_33848)
  );
  InMux inmux_8_2_33814_33841 (
    .I(net_33814),
    .O(net_33841)
  );
  InMux inmux_8_2_33814_33855 (
    .I(net_33814),
    .O(net_33855)
  );
  InMux inmux_8_2_33814_33858 (
    .I(net_33814),
    .O(net_33858)
  );
  InMux inmux_8_2_33814_33867 (
    .I(net_33814),
    .O(net_33867)
  );
  InMux inmux_8_2_33815_33830 (
    .I(net_33815),
    .O(net_33830)
  );
  InMux inmux_8_2_33815_33842 (
    .I(net_33815),
    .O(net_33842)
  );
  InMux inmux_8_2_33815_33847 (
    .I(net_33815),
    .O(net_33847)
  );
  InMux inmux_8_2_33815_33854 (
    .I(net_33815),
    .O(net_33854)
  );
  InMux inmux_8_2_33815_33859 (
    .I(net_33815),
    .O(net_33859)
  );
  InMux inmux_8_2_33815_33866 (
    .I(net_33815),
    .O(net_33866)
  );
  CEMux inmux_8_2_33816_33868 (
    .I(net_33816),
    .O(net_33868)
  );
  InMux inmux_8_2_33817_33840 (
    .I(net_33817),
    .O(net_33840)
  );
  InMux inmux_8_2_33817_33852 (
    .I(net_33817),
    .O(net_33852)
  );
  InMux inmux_8_2_33817_33861 (
    .I(net_33817),
    .O(net_33861)
  );
  InMux inmux_8_2_33817_33864 (
    .I(net_33817),
    .O(net_33864)
  );
  ClkMux inmux_8_2_5_33869 (
    .I(net_5),
    .O(net_33869)
  );
  IoInMux inmux_8_31_37376_37363 (
    .I(net_37376),
    .O(net_37363)
  );
  CEMux inmux_8_31_37382_37366 (
    .I(net_37382),
    .O(net_37366)
  );
  ClkMux inmux_8_31_5_37367 (
    .I(net_5),
    .O(net_37367)
  );
  ClkMux inmux_8_31_5_37368 (
    .I(net_5),
    .O(net_37368)
  );
  InMux inmux_8_3_33912_33952 (
    .I(net_33912),
    .O(net_33952)
  );
  InMux inmux_8_3_33912_33988 (
    .I(net_33912),
    .O(net_33988)
  );
  CEMux inmux_8_3_33914_33991 (
    .I(net_33914),
    .O(net_33991)
  );
  InMux inmux_8_3_33916_33954 (
    .I(net_33916),
    .O(net_33954)
  );
  InMux inmux_8_3_33926_33987 (
    .I(net_33926),
    .O(net_33987)
  );
  InMux inmux_8_3_33929_33970 (
    .I(net_33929),
    .O(net_33970)
  );
  InMux inmux_8_3_33929_33977 (
    .I(net_33929),
    .O(net_33977)
  );
  InMux inmux_8_3_33929_33984 (
    .I(net_33929),
    .O(net_33984)
  );
  InMux inmux_8_3_33932_33971 (
    .I(net_33932),
    .O(net_33971)
  );
  InMux inmux_8_3_33932_33978 (
    .I(net_33932),
    .O(net_33978)
  );
  InMux inmux_8_3_33932_33983 (
    .I(net_33932),
    .O(net_33983)
  );
  InMux inmux_8_3_33938_33972 (
    .I(net_33938),
    .O(net_33972)
  );
  InMux inmux_8_3_33938_33975 (
    .I(net_33938),
    .O(net_33975)
  );
  InMux inmux_8_3_33938_33982 (
    .I(net_33938),
    .O(net_33982)
  );
  InMux inmux_8_3_33941_33969 (
    .I(net_33941),
    .O(net_33969)
  );
  InMux inmux_8_3_33941_33976 (
    .I(net_33941),
    .O(net_33976)
  );
  InMux inmux_8_3_33941_33981 (
    .I(net_33941),
    .O(net_33981)
  );
  ClkMux inmux_8_3_5_33992 (
    .I(net_5),
    .O(net_33992)
  );
  InMux inmux_9_10_38610_38644 (
    .I(net_38610),
    .O(net_38644)
  );
  InMux inmux_9_10_38610_38649 (
    .I(net_38610),
    .O(net_38649)
  );
  InMux inmux_9_10_38610_38675 (
    .I(net_38610),
    .O(net_38675)
  );
  CEMux inmux_9_10_38622_38683 (
    .I(net_38622),
    .O(net_38683)
  );
  InMux inmux_9_10_38627_38645 (
    .I(net_38627),
    .O(net_38645)
  );
  InMux inmux_9_10_38627_38674 (
    .I(net_38627),
    .O(net_38674)
  );
  InMux inmux_9_10_38630_38643 (
    .I(net_38630),
    .O(net_38643)
  );
  InMux inmux_9_10_38630_38676 (
    .I(net_38630),
    .O(net_38676)
  );
  InMux inmux_9_10_38632_38681 (
    .I(net_38632),
    .O(net_38681)
  );
  InMux inmux_9_10_38635_38646 (
    .I(net_38635),
    .O(net_38646)
  );
  InMux inmux_9_10_38635_38661 (
    .I(net_38635),
    .O(net_38661)
  );
  InMux inmux_9_10_38635_38673 (
    .I(net_38635),
    .O(net_38673)
  );
  ClkMux inmux_9_10_5_38684 (
    .I(net_5),
    .O(net_38684)
  );
  InMux inmux_9_11_38745_38793 (
    .I(net_38745),
    .O(net_38793)
  );
  ClkMux inmux_9_11_5_38807 (
    .I(net_5),
    .O(net_38807)
  );
  CEMux inmux_9_11_6_38806 (
    .I(net_6),
    .O(net_38806)
  );
  InMux inmux_9_12_38864_38891 (
    .I(net_38864),
    .O(net_38891)
  );
  CEMux inmux_9_12_38868_38929 (
    .I(net_38868),
    .O(net_38929)
  );
  ClkMux inmux_9_12_5_38930 (
    .I(net_5),
    .O(net_38930)
  );
  InMux inmux_9_18_39609_39629 (
    .I(net_39609),
    .O(net_39629)
  );
  InMux inmux_9_18_39610_39654 (
    .I(net_39610),
    .O(net_39654)
  );
  ClkMux inmux_9_18_5_39668 (
    .I(net_5),
    .O(net_39668)
  );
  CEMux inmux_9_18_6_39667 (
    .I(net_6),
    .O(net_39667)
  );
  InMux inmux_9_27_40696_40770 (
    .I(net_40696),
    .O(net_40770)
  );
  CEMux inmux_9_27_40706_40774 (
    .I(net_40706),
    .O(net_40774)
  );
  InMux inmux_9_27_40715_40761 (
    .I(net_40715),
    .O(net_40761)
  );
  InMux inmux_9_27_40715_40771 (
    .I(net_40715),
    .O(net_40771)
  );
  InMux inmux_9_27_40718_40736 (
    .I(net_40718),
    .O(net_40736)
  );
  InMux inmux_9_27_40719_40734 (
    .I(net_40719),
    .O(net_40734)
  );
  InMux inmux_9_27_40721_40760 (
    .I(net_40721),
    .O(net_40760)
  );
  ClkMux inmux_9_27_5_40775 (
    .I(net_5),
    .O(net_40775)
  );
  InMux inmux_9_28_40818_40865 (
    .I(net_40818),
    .O(net_40865)
  );
  InMux inmux_9_28_40820_40887 (
    .I(net_40820),
    .O(net_40887)
  );
  InMux inmux_9_28_40823_40859 (
    .I(net_40823),
    .O(net_40859)
  );
  InMux inmux_9_28_40825_40890 (
    .I(net_40825),
    .O(net_40890)
  );
  InMux inmux_9_28_40826_40866 (
    .I(net_40826),
    .O(net_40866)
  );
  InMux inmux_9_28_40828_40857 (
    .I(net_40828),
    .O(net_40857)
  );
  InMux inmux_9_28_40831_40889 (
    .I(net_40831),
    .O(net_40889)
  );
  InMux inmux_9_28_40833_40882 (
    .I(net_40833),
    .O(net_40882)
  );
  CEMux inmux_9_28_40836_40897 (
    .I(net_40836),
    .O(net_40897)
  );
  InMux inmux_9_28_40837_40888 (
    .I(net_40837),
    .O(net_40888)
  );
  InMux inmux_9_28_40839_40864 (
    .I(net_40839),
    .O(net_40864)
  );
  ClkMux inmux_9_28_5_40898 (
    .I(net_5),
    .O(net_40898)
  );
  InMux inmux_9_29_40941_40993 (
    .I(net_40941),
    .O(net_40993)
  );
  InMux inmux_9_29_40950_40995 (
    .I(net_40950),
    .O(net_40995)
  );
  InMux inmux_9_29_40957_40976 (
    .I(net_40957),
    .O(net_40976)
  );
  InMux inmux_9_29_40960_40977 (
    .I(net_40960),
    .O(net_40977)
  );
  InMux inmux_9_29_40960_41006 (
    .I(net_40960),
    .O(net_41006)
  );
  InMux inmux_9_29_40961_40974 (
    .I(net_40961),
    .O(net_40974)
  );
  InMux inmux_9_29_40961_41005 (
    .I(net_40961),
    .O(net_41005)
  );
  InMux inmux_9_29_40962_40975 (
    .I(net_40962),
    .O(net_40975)
  );
  InMux inmux_9_29_40965_41004 (
    .I(net_40965),
    .O(net_41004)
  );
  InMux inmux_9_29_40970_41007 (
    .I(net_40970),
    .O(net_41007)
  );
  InMux inmux_9_2_37621_37678 (
    .I(net_37621),
    .O(net_37678)
  );
  InMux inmux_9_2_37622_37679 (
    .I(net_37622),
    .O(net_37679)
  );
  InMux inmux_9_2_37623_37690 (
    .I(net_37623),
    .O(net_37690)
  );
  InMux inmux_9_2_37624_37689 (
    .I(net_37624),
    .O(net_37689)
  );
  InMux inmux_9_2_37627_37692 (
    .I(net_37627),
    .O(net_37692)
  );
  CEMux inmux_9_2_37631_37699 (
    .I(net_37631),
    .O(net_37699)
  );
  InMux inmux_9_2_37632_37680 (
    .I(net_37632),
    .O(net_37680)
  );
  InMux inmux_9_2_37633_37662 (
    .I(net_37633),
    .O(net_37662)
  );
  InMux inmux_9_2_37635_37674 (
    .I(net_37635),
    .O(net_37674)
  );
  InMux inmux_9_2_37637_37654 (
    .I(net_37637),
    .O(net_37654)
  );
  InMux inmux_9_2_37638_37691 (
    .I(net_37638),
    .O(net_37691)
  );
  InMux inmux_9_2_37639_37659 (
    .I(net_37639),
    .O(net_37659)
  );
  InMux inmux_9_2_37639_37661 (
    .I(net_37639),
    .O(net_37661)
  );
  InMux inmux_9_2_37640_37653 (
    .I(net_37640),
    .O(net_37653)
  );
  InMux inmux_9_2_37640_37667 (
    .I(net_37640),
    .O(net_37667)
  );
  InMux inmux_9_2_37642_37655 (
    .I(net_37642),
    .O(net_37655)
  );
  InMux inmux_9_2_37642_37698 (
    .I(net_37642),
    .O(net_37698)
  );
  InMux inmux_9_2_37643_37656 (
    .I(net_37643),
    .O(net_37656)
  );
  InMux inmux_9_2_37646_37668 (
    .I(net_37646),
    .O(net_37668)
  );
  InMux inmux_9_2_37647_37684 (
    .I(net_37647),
    .O(net_37684)
  );
  InMux inmux_9_2_37647_37696 (
    .I(net_37647),
    .O(net_37696)
  );
  InMux inmux_9_2_37648_37673 (
    .I(net_37648),
    .O(net_37673)
  );
  InMux inmux_9_2_37649_37677 (
    .I(net_37649),
    .O(net_37677)
  );
  InMux inmux_9_2_37650_37666 (
    .I(net_37650),
    .O(net_37666)
  );
  InMux inmux_9_2_37651_37665 (
    .I(net_37651),
    .O(net_37665)
  );
  ClkMux inmux_9_2_5_37700 (
    .I(net_5),
    .O(net_37700)
  );
  InMux inmux_9_30_41064_41140 (
    .I(net_41064),
    .O(net_41140)
  );
  InMux inmux_9_30_41068_41142 (
    .I(net_41068),
    .O(net_41142)
  );
  InMux inmux_9_30_41072_41098 (
    .I(net_41072),
    .O(net_41098)
  );
  InMux inmux_9_30_41072_41112 (
    .I(net_41072),
    .O(net_41112)
  );
  InMux inmux_9_30_41072_41139 (
    .I(net_41072),
    .O(net_41139)
  );
  InMux inmux_9_30_41077_41099 (
    .I(net_41077),
    .O(net_41099)
  );
  InMux inmux_9_30_41077_41109 (
    .I(net_41077),
    .O(net_41109)
  );
  CEMux inmux_9_30_41082_41143 (
    .I(net_41082),
    .O(net_41143)
  );
  InMux inmux_9_30_41083_41100 (
    .I(net_41083),
    .O(net_41100)
  );
  InMux inmux_9_30_41083_41110 (
    .I(net_41083),
    .O(net_41110)
  );
  InMux inmux_9_30_41084_41097 (
    .I(net_41084),
    .O(net_41097)
  );
  InMux inmux_9_30_41084_41111 (
    .I(net_41084),
    .O(net_41111)
  );
  InMux inmux_9_30_41094_41127 (
    .I(net_41094),
    .O(net_41127)
  );
  ClkMux inmux_9_30_5_41144 (
    .I(net_5),
    .O(net_41144)
  );
  InMux inmux_9_3_37748_37791 (
    .I(net_37748),
    .O(net_37791)
  );
  InMux inmux_9_3_37748_37806 (
    .I(net_37748),
    .O(net_37806)
  );
  InMux inmux_9_3_37748_37813 (
    .I(net_37748),
    .O(net_37813)
  );
  InMux inmux_9_3_37748_37818 (
    .I(net_37748),
    .O(net_37818)
  );
  InMux inmux_9_3_37749_37783 (
    .I(net_37749),
    .O(net_37783)
  );
  InMux inmux_9_3_37749_37800 (
    .I(net_37749),
    .O(net_37800)
  );
  InMux inmux_9_3_37752_37790 (
    .I(net_37752),
    .O(net_37790)
  );
  InMux inmux_9_3_37752_37807 (
    .I(net_37752),
    .O(net_37807)
  );
  InMux inmux_9_3_37752_37812 (
    .I(net_37752),
    .O(net_37812)
  );
  InMux inmux_9_3_37752_37819 (
    .I(net_37752),
    .O(net_37819)
  );
  CEMux inmux_9_3_37754_37822 (
    .I(net_37754),
    .O(net_37822)
  );
  InMux inmux_9_3_37755_37808 (
    .I(net_37755),
    .O(net_37808)
  );
  InMux inmux_9_3_37756_37797 (
    .I(net_37756),
    .O(net_37797)
  );
  InMux inmux_9_3_37757_37784 (
    .I(net_37757),
    .O(net_37784)
  );
  InMux inmux_9_3_37759_37776 (
    .I(net_37759),
    .O(net_37776)
  );
  InMux inmux_9_3_37760_37777 (
    .I(net_37760),
    .O(net_37777)
  );
  InMux inmux_9_3_37760_37794 (
    .I(net_37760),
    .O(net_37794)
  );
  InMux inmux_9_3_37763_37778 (
    .I(net_37763),
    .O(net_37778)
  );
  InMux inmux_9_3_37763_37785 (
    .I(net_37763),
    .O(net_37785)
  );
  InMux inmux_9_3_37763_37788 (
    .I(net_37763),
    .O(net_37788)
  );
  InMux inmux_9_3_37763_37795 (
    .I(net_37763),
    .O(net_37795)
  );
  InMux inmux_9_3_37763_37821 (
    .I(net_37763),
    .O(net_37821)
  );
  InMux inmux_9_3_37764_37803 (
    .I(net_37764),
    .O(net_37803)
  );
  InMux inmux_9_3_37766_37801 (
    .I(net_37766),
    .O(net_37801)
  );
  InMux inmux_9_3_37768_37809 (
    .I(net_37768),
    .O(net_37809)
  );
  InMux inmux_9_3_37768_37814 (
    .I(net_37768),
    .O(net_37814)
  );
  InMux inmux_9_3_37769_37779 (
    .I(net_37769),
    .O(net_37779)
  );
  InMux inmux_9_3_37769_37789 (
    .I(net_37769),
    .O(net_37789)
  );
  InMux inmux_9_3_37769_37796 (
    .I(net_37769),
    .O(net_37796)
  );
  InMux inmux_9_3_37769_37815 (
    .I(net_37769),
    .O(net_37815)
  );
  InMux inmux_9_3_37769_37820 (
    .I(net_37769),
    .O(net_37820)
  );
  InMux inmux_9_3_37770_37802 (
    .I(net_37770),
    .O(net_37802)
  );
  ClkMux inmux_9_3_5_37823 (
    .I(net_5),
    .O(net_37823)
  );
  InMux inmux_9_4_37866_37901 (
    .I(net_37866),
    .O(net_37901)
  );
  InMux inmux_9_4_37869_37905 (
    .I(net_37869),
    .O(net_37905)
  );
  InMux inmux_9_4_37869_37931 (
    .I(net_37869),
    .O(net_37931)
  );
  CEMux inmux_9_4_37877_37945 (
    .I(net_37877),
    .O(net_37945)
  );
  InMux inmux_9_4_37883_37929 (
    .I(net_37883),
    .O(net_37929)
  );
  InMux inmux_9_4_37895_37899 (
    .I(net_37895),
    .O(net_37899)
  );
  InMux inmux_9_4_37895_37930 (
    .I(net_37895),
    .O(net_37930)
  );
  ClkMux inmux_9_4_5_37946 (
    .I(net_5),
    .O(net_37946)
  );
  CEMux inmux_9_5_38000_38068 (
    .I(net_38000),
    .O(net_38068)
  );
  InMux inmux_9_5_38014_38041 (
    .I(net_38014),
    .O(net_38041)
  );
  ClkMux inmux_9_5_5_38069 (
    .I(net_5),
    .O(net_38069)
  );
  InMux inmux_9_8_38364_38417 (
    .I(net_38364),
    .O(net_38417)
  );
  InMux inmux_9_8_38367_38393 (
    .I(net_38367),
    .O(net_38393)
  );
  InMux inmux_9_8_38373_38398 (
    .I(net_38373),
    .O(net_38398)
  );
  InMux inmux_9_8_38376_38429 (
    .I(net_38376),
    .O(net_38429)
  );
  InMux inmux_9_8_38380_38434 (
    .I(net_38380),
    .O(net_38434)
  );
  InMux inmux_9_8_38382_38411 (
    .I(net_38382),
    .O(net_38411)
  );
  InMux inmux_9_8_38383_38405 (
    .I(net_38383),
    .O(net_38405)
  );
  InMux inmux_9_8_38386_38423 (
    .I(net_38386),
    .O(net_38423)
  );
  InMux inmux_9_8_38396_38406 (
    .I(net_38396),
    .O(net_38406)
  );
  InMux inmux_9_8_38402_38412 (
    .I(net_38402),
    .O(net_38412)
  );
  InMux inmux_9_8_38408_38418 (
    .I(net_38408),
    .O(net_38418)
  );
  InMux inmux_9_8_38414_38424 (
    .I(net_38414),
    .O(net_38424)
  );
  InMux inmux_9_8_38420_38430 (
    .I(net_38420),
    .O(net_38430)
  );
  InMux inmux_9_8_38426_38436 (
    .I(net_38426),
    .O(net_38436)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_42481),
    .in2(net_42482_cascademuxed),
    .in3(gnd),
    .lcout(net_38565),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42593_cascademuxed),
    .in3(gnd),
    .lcout(net_38686),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_42597),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38687),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42637),
    .clk(net_42638),
    .in0(net_42603),
    .in1(gnd),
    .in2(net_42605_cascademuxed),
    .in3(net_42606),
    .lcout(net_38688),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42618),
    .lcout(net_38690),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_12_0 (
    .carryin(t109),
    .carryout(net_42713),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_42715),
    .in2(net_42716_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_12_1 (
    .carryin(net_42713),
    .carryout(net_42719),
    .ce(net_42760),
    .clk(net_42761),
    .in0(gnd),
    .in1(net_42721),
    .in2(net_42722_cascademuxed),
    .in3(net_42723),
    .lcout(net_38810),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_12_2 (
    .carryin(net_42719),
    .carryout(net_42725),
    .ce(net_42760),
    .clk(net_42761),
    .in0(gnd),
    .in1(net_42727),
    .in2(net_42728_cascademuxed),
    .in3(net_42729),
    .lcout(net_38811),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_12_3 (
    .carryin(net_42725),
    .carryout(net_42731),
    .ce(net_42760),
    .clk(net_42761),
    .in0(gnd),
    .in1(net_42733),
    .in2(net_42734_cascademuxed),
    .in3(net_42735),
    .lcout(net_38812),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_12_4 (
    .carryin(net_42731),
    .carryout(net_42737),
    .ce(net_42760),
    .clk(net_42761),
    .in0(gnd),
    .in1(net_42739),
    .in2(net_42740_cascademuxed),
    .in3(net_42741),
    .lcout(net_38813),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_12_5 (
    .carryin(net_42737),
    .carryout(net_42743),
    .ce(net_42760),
    .clk(net_42761),
    .in0(gnd),
    .in1(net_42745),
    .in2(net_42746_cascademuxed),
    .in3(net_42747),
    .lcout(net_38814),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_12_6 (
    .carryin(net_42743),
    .carryout(net_42749),
    .ce(net_42760),
    .clk(net_42761),
    .in0(gnd),
    .in1(net_42751),
    .in2(net_42752_cascademuxed),
    .in3(net_42753),
    .lcout(net_38815),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_12_7 (
    .carryin(net_42749),
    .carryout(net_42755),
    .ce(net_42760),
    .clk(net_42761),
    .in0(gnd),
    .in1(net_42757),
    .in2(net_42758_cascademuxed),
    .in3(net_42759),
    .lcout(net_38816),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_0 (
    .carryin(net_42799),
    .carryout(net_42836),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(net_42838),
    .in2(net_42839_cascademuxed),
    .in3(net_42840),
    .lcout(net_38932),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_1 (
    .carryin(net_42836),
    .carryout(net_42842),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(net_42844),
    .in2(net_42845_cascademuxed),
    .in3(net_42846),
    .lcout(net_38933),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_2 (
    .carryin(net_42842),
    .carryout(net_42848),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(net_42850),
    .in2(net_42851_cascademuxed),
    .in3(net_42852),
    .lcout(net_38934),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_3 (
    .carryin(net_42848),
    .carryout(net_42854),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(net_42856),
    .in2(net_42857_cascademuxed),
    .in3(net_42858),
    .lcout(net_38935),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_4 (
    .carryin(net_42854),
    .carryout(net_42860),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(net_42862),
    .in2(net_42863_cascademuxed),
    .in3(net_42864),
    .lcout(net_38936),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_5 (
    .carryin(net_42860),
    .carryout(net_42866),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(net_42868),
    .in2(net_42869_cascademuxed),
    .in3(net_42870),
    .lcout(net_38937),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_6 (
    .carryin(net_42866),
    .carryout(net_42872),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(net_42874),
    .in2(net_42875_cascademuxed),
    .in3(net_42876),
    .lcout(net_38938),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42883),
    .clk(net_42884),
    .in0(gnd),
    .in1(net_42880),
    .in2(net_42881_cascademuxed),
    .in3(net_42882),
    .lcout(net_38939),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42962_cascademuxed),
    .in3(gnd),
    .lcout(net_39055),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42969),
    .lcout(net_39056),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42974_cascademuxed),
    .in3(gnd),
    .lcout(net_39057),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42981),
    .lcout(net_39058),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(net_42984),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39059),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42992_cascademuxed),
    .in3(gnd),
    .lcout(net_39060),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_42998_cascademuxed),
    .in3(gnd),
    .lcout(net_39061),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43006),
    .clk(net_43007),
    .in0(gnd),
    .in1(net_43003),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39062),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43085_cascademuxed),
    .in3(gnd),
    .lcout(net_39178),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_10_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_43129),
    .clk(net_43130),
    .in0(gnd),
    .in1(net_43096),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_39180),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43109_cascademuxed),
    .in3(gnd),
    .lcout(net_39182),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_17_0 (
    .carryin(t113),
    .carryout(t115),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43331_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_17_1 (
    .carryin(t115),
    .carryout(net_43334),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_43336),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_2 (
    .carryin(net_43334),
    .carryout(net_43340),
    .ce(),
    .clk(net_43376),
    .in0(gnd),
    .in1(net_43342),
    .in2(gnd),
    .in3(net_43344),
    .lcout(net_39426),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_3 (
    .carryin(net_43340),
    .carryout(net_43346),
    .ce(),
    .clk(net_43376),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43349_cascademuxed),
    .in3(net_43350),
    .lcout(net_39427),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_4 (
    .carryin(net_43346),
    .carryout(net_43352),
    .ce(),
    .clk(net_43376),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43355_cascademuxed),
    .in3(net_43356),
    .lcout(net_39428),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_5 (
    .carryin(net_43352),
    .carryout(net_43358),
    .ce(),
    .clk(net_43376),
    .in0(gnd),
    .in1(net_43360),
    .in2(gnd),
    .in3(net_43362),
    .lcout(net_39429),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_6 (
    .carryin(net_43358),
    .carryout(net_43364),
    .ce(),
    .clk(net_43376),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43367_cascademuxed),
    .in3(net_43368),
    .lcout(net_39430),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_17_7 (
    .carryin(net_43364),
    .carryout(net_43370),
    .ce(),
    .clk(net_43376),
    .in0(gnd),
    .in1(net_43372),
    .in2(gnd),
    .in3(net_43374),
    .lcout(net_39431),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_0 (
    .carryin(net_43414),
    .carryout(net_43451),
    .ce(),
    .clk(net_43499),
    .in0(gnd),
    .in1(net_43453),
    .in2(gnd),
    .in3(net_43455),
    .lcout(net_39547),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_1 (
    .carryin(net_43451),
    .carryout(net_43457),
    .ce(),
    .clk(net_43499),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43460_cascademuxed),
    .in3(net_43461),
    .lcout(net_39548),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_2 (
    .carryin(net_43457),
    .carryout(net_43463),
    .ce(),
    .clk(net_43499),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43466_cascademuxed),
    .in3(net_43467),
    .lcout(net_39549),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_3 (
    .carryin(net_43463),
    .carryout(net_43469),
    .ce(),
    .clk(net_43499),
    .in0(gnd),
    .in1(net_43471),
    .in2(gnd),
    .in3(net_43473),
    .lcout(net_39550),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_4 (
    .carryin(net_43469),
    .carryout(net_43475),
    .ce(),
    .clk(net_43499),
    .in0(gnd),
    .in1(net_43477),
    .in2(gnd),
    .in3(net_43479),
    .lcout(net_39551),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_5 (
    .carryin(net_43475),
    .carryout(net_43481),
    .ce(),
    .clk(net_43499),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43484_cascademuxed),
    .in3(net_43485),
    .lcout(net_39552),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_6 (
    .carryin(net_43481),
    .carryout(net_43487),
    .ce(),
    .clk(net_43499),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43490_cascademuxed),
    .in3(net_43491),
    .lcout(net_39553),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_18_7 (
    .carryin(net_43487),
    .carryout(net_43493),
    .ce(),
    .clk(net_43499),
    .in0(gnd),
    .in1(net_43495),
    .in2(gnd),
    .in3(net_43497),
    .lcout(net_39554),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_0 (
    .carryin(net_43537),
    .carryout(net_43574),
    .ce(),
    .clk(net_43622),
    .in0(gnd),
    .in1(net_43576),
    .in2(gnd),
    .in3(net_43578),
    .lcout(net_39670),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_1 (
    .carryin(net_43574),
    .carryout(net_43580),
    .ce(),
    .clk(net_43622),
    .in0(gnd),
    .in1(net_43582),
    .in2(gnd),
    .in3(net_43584),
    .lcout(net_39671),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_2 (
    .carryin(net_43580),
    .carryout(net_43586),
    .ce(),
    .clk(net_43622),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43589_cascademuxed),
    .in3(net_43590),
    .lcout(net_39672),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_3 (
    .carryin(net_43586),
    .carryout(net_43592),
    .ce(),
    .clk(net_43622),
    .in0(gnd),
    .in1(net_43594),
    .in2(gnd),
    .in3(net_43596),
    .lcout(net_39673),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_4 (
    .carryin(net_43592),
    .carryout(net_43598),
    .ce(),
    .clk(net_43622),
    .in0(gnd),
    .in1(net_43600),
    .in2(gnd),
    .in3(net_43602),
    .lcout(net_39674),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_5 (
    .carryin(net_43598),
    .carryout(net_43604),
    .ce(),
    .clk(net_43622),
    .in0(gnd),
    .in1(net_43606),
    .in2(gnd),
    .in3(net_43608),
    .lcout(net_39675),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_6 (
    .carryin(net_43604),
    .carryout(net_43610),
    .ce(),
    .clk(net_43622),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43613_cascademuxed),
    .in3(net_43614),
    .lcout(net_39676),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_19_7 (
    .carryin(net_43610),
    .carryout(net_43616),
    .ce(),
    .clk(net_43622),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43619_cascademuxed),
    .in3(net_43620),
    .lcout(net_39677),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_1_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_20_0 (
    .carryin(net_43660),
    .carryout(net_43697),
    .ce(),
    .clk(net_43745),
    .in0(gnd),
    .in1(net_43699),
    .in2(gnd),
    .in3(net_43701),
    .lcout(net_39793),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_20_1 (
    .carryin(net_43697),
    .carryout(net_43703),
    .ce(),
    .clk(net_43745),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43706_cascademuxed),
    .in3(net_43707),
    .lcout(net_39794),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_20_2 (
    .carryin(net_43703),
    .carryout(net_43709),
    .ce(),
    .clk(net_43745),
    .in0(gnd),
    .in1(net_43711),
    .in2(gnd),
    .in3(net_43713),
    .lcout(net_39795),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_20_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_43745),
    .in0(gnd),
    .in1(gnd),
    .in2(net_43718_cascademuxed),
    .in3(net_43719),
    .lcout(net_39796),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_26_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44448),
    .in1(gnd),
    .in2(gnd),
    .in3(net_44451),
    .lcout(net_40533),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_26_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44482),
    .clk(net_44483),
    .in0(net_44478),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_40538),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_27_0 (
    .carryin(t120),
    .carryout(t122),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_44561_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_27_1 (
    .carryin(t122),
    .carryout(net_44564),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_44567_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_27_2 (
    .carryin(net_44564),
    .carryout(net_44570),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_44572),
    .in2(gnd),
    .in3(net_44574),
    .lcout(net_40656),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_27_3 (
    .carryin(net_44570),
    .carryout(net_44576),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_44579_cascademuxed),
    .in3(net_44580),
    .lcout(net_40657),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_27_4 (
    .carryin(net_44576),
    .carryout(net_44582),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_44584),
    .in2(gnd),
    .in3(net_44586),
    .lcout(net_40658),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_27_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_44590),
    .in2(gnd),
    .in3(net_44592),
    .lcout(net_40659),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_27_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44605),
    .clk(net_44606),
    .in0(net_44595),
    .in1(net_44596),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_40660),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_27_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44605),
    .clk(net_44606),
    .in0(net_44601),
    .in1(gnd),
    .in2(gnd),
    .in3(net_44604),
    .lcout(net_40661),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_28_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44694),
    .in1(net_44695),
    .in2(net_44696_cascademuxed),
    .in3(net_44697),
    .lcout(net_40779),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000001000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_28_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44728),
    .clk(net_44729),
    .in0(gnd),
    .in1(net_44701),
    .in2(net_44702_cascademuxed),
    .in3(net_44703),
    .lcout(net_40780),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_28_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44712),
    .in1(net_44713),
    .in2(net_44714_cascademuxed),
    .in3(net_44715),
    .lcout(net_40782),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_28_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44728),
    .clk(net_44729),
    .in0(gnd),
    .in1(gnd),
    .in2(net_44726_cascademuxed),
    .in3(net_44727),
    .lcout(net_40784),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001101010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_29_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44851),
    .clk(net_44852),
    .in0(net_44805),
    .in1(net_44806),
    .in2(net_44807_cascademuxed),
    .in3(net_44808),
    .lcout(net_40900),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_10_29_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44817),
    .in1(net_44818),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_40902),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_29_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44823),
    .in1(net_44824),
    .in2(net_44825_cascademuxed),
    .in3(net_44826),
    .lcout(net_40903),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100000110000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_29_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44851),
    .clk(net_44852),
    .in0(net_44835),
    .in1(net_44836),
    .in2(net_44837_cascademuxed),
    .in3(net_44838),
    .lcout(net_40905),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_29_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44841),
    .in1(net_44842),
    .in2(net_44843_cascademuxed),
    .in3(net_44844),
    .lcout(net_40906),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111000010000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_29_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44847),
    .in1(net_44848),
    .in2(net_44849_cascademuxed),
    .in3(net_44850),
    .lcout(net_40907),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_2_0 (
    .carryin(t81),
    .carryout(t83),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_41485),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_2_1 (
    .carryin(t83),
    .carryout(net_41489),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_41491),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_2_2 (
    .carryin(net_41489),
    .carryout(net_41495),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_41497),
    .in2(gnd),
    .in3(net_41499),
    .lcout(net_37545),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_2_3 (
    .carryin(net_41495),
    .carryout(net_41501),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41504_cascademuxed),
    .in3(net_41505),
    .lcout(net_37546),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_2_4 (
    .carryin(net_41501),
    .carryout(net_41507),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_41509),
    .in2(gnd),
    .in3(net_41511),
    .lcout(net_37547),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_41515),
    .in2(gnd),
    .in3(net_41517),
    .lcout(net_37548),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41530),
    .clk(net_41531),
    .in0(net_41520),
    .in1(gnd),
    .in2(net_41522_cascademuxed),
    .in3(gnd),
    .lcout(net_37549),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41530),
    .clk(net_41531),
    .in0(net_41526),
    .in1(gnd),
    .in2(gnd),
    .in3(net_41529),
    .lcout(net_37550),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_10_30_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_44929),
    .in2(net_44930_cascademuxed),
    .in3(gnd),
    .lcout(net_41023),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0111011000010001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_30_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44940),
    .in1(net_44941),
    .in2(net_44942_cascademuxed),
    .in3(net_44943),
    .lcout(net_41025),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011111010101010),
    .SEQ_MODE(4'b1000)
  ) lc40_10_30_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44974),
    .clk(net_44975),
    .in0(net_44946),
    .in1(net_44947),
    .in2(net_44948_cascademuxed),
    .in3(net_44949),
    .lcout(net_41026),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111011011110),
    .SEQ_MODE(4'b1000)
  ) lc40_10_30_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_44974),
    .clk(net_44975),
    .in0(net_44952),
    .in1(net_44953),
    .in2(net_44954_cascademuxed),
    .in3(net_44955),
    .lcout(net_41027),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101101000011010),
    .SEQ_MODE(4'b0000)
  ) lc40_10_30_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44964),
    .in1(net_44965),
    .in2(net_44966_cascademuxed),
    .in3(net_44967),
    .lcout(net_41029),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110000111110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_30_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_44970),
    .in1(net_44971),
    .in2(net_44972_cascademuxed),
    .in3(net_44973),
    .lcout(net_41030),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41653),
    .clk(net_41654),
    .in0(net_41619),
    .in1(gnd),
    .in2(net_41621_cascademuxed),
    .in3(gnd),
    .lcout(net_37704),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41653),
    .clk(net_41654),
    .in0(gnd),
    .in1(net_41626),
    .in2(gnd),
    .in3(net_41628),
    .lcout(net_37705),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41653),
    .clk(net_41654),
    .in0(net_41631),
    .in1(gnd),
    .in2(net_41633_cascademuxed),
    .in3(gnd),
    .lcout(net_37706),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000101000),
    .SEQ_MODE(4'b1000)
  ) lc40_10_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41653),
    .clk(net_41654),
    .in0(net_41643),
    .in1(net_41644),
    .in2(net_41645_cascademuxed),
    .in3(gnd),
    .lcout(net_37708),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_10_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_41651_cascademuxed),
    .in3(net_41652),
    .lcout(net_37709),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000010),
    .SEQ_MODE(4'b0000)
  ) lc40_10_7_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_42129),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42132),
    .lcout(net_38199),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000010111111),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42268),
    .clk(net_42269),
    .in0(net_42222),
    .in1(net_42223),
    .in2(net_42224_cascademuxed),
    .in3(net_42225),
    .lcout(net_38317),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_10_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_42228),
    .in1(net_42229),
    .in2(net_42230_cascademuxed),
    .in3(net_42231),
    .lcout(net_38318),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_8_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_42237),
    .lcout(net_38319),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001101010011),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42268),
    .clk(net_42269),
    .in0(net_42240),
    .in1(net_42241),
    .in2(net_42242_cascademuxed),
    .in3(net_42243),
    .lcout(net_38320),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_42246),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38321),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_10_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_42258),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_38323),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001100011011),
    .SEQ_MODE(4'b1000)
  ) lc40_10_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_42268),
    .clk(net_42269),
    .in0(net_42264),
    .in1(net_42265),
    .in2(net_42266_cascademuxed),
    .in3(net_42267),
    .lcout(net_38324),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100110000001100),
    .SEQ_MODE(4'b0000)
  ) lc40_11_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46299),
    .in1(net_46300),
    .in2(net_46301_cascademuxed),
    .in3(net_46302),
    .lcout(net_42394),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46317),
    .in1(gnd),
    .in2(net_46319_cascademuxed),
    .in3(gnd),
    .lcout(net_42397),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46345),
    .clk(net_46346),
    .in0(gnd),
    .in1(net_46324),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42398),
    .ltout(),
    .sr(net_46347)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46329),
    .in1(gnd),
    .in2(net_46331_cascademuxed),
    .in3(gnd),
    .lcout(net_42399),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010101),
    .SEQ_MODE(4'b0000)
  ) lc40_11_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46336),
    .in2(net_46337_cascademuxed),
    .in3(net_46338),
    .lcout(net_42400),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46341),
    .in1(net_46342),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42401),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46468),
    .clk(net_46469),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46436_cascademuxed),
    .in3(gnd),
    .lcout(net_42519),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46468),
    .clk(net_46469),
    .in0(net_46464),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42524),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001110100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46551),
    .in1(net_46552),
    .in2(net_46553_cascademuxed),
    .in3(net_46554),
    .lcout(net_42641),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46591),
    .clk(net_46592),
    .in0(net_46557),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42642),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111101110111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46563),
    .in1(net_46564),
    .in2(net_46565_cascademuxed),
    .in3(net_46566),
    .lcout(net_42643),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46569),
    .in1(net_46570),
    .in2(net_46571_cascademuxed),
    .in3(net_46572),
    .lcout(net_42644),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46581),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42646),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46591),
    .clk(net_46592),
    .in0(gnd),
    .in1(net_46588),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42647),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101001101011111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46668),
    .in1(net_46669),
    .in2(net_46670_cascademuxed),
    .in3(net_46671),
    .lcout(net_42763),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100011101110111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46674),
    .in1(net_46675),
    .in2(net_46676_cascademuxed),
    .in3(net_46677),
    .lcout(net_42764),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010110111111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46680),
    .in1(net_46681),
    .in2(net_46682_cascademuxed),
    .in3(net_46683),
    .lcout(net_42765),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46688_cascademuxed),
    .in3(gnd),
    .lcout(net_42766),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011111110111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46692),
    .in1(net_46693),
    .in2(net_46694_cascademuxed),
    .in3(net_46695),
    .lcout(net_42767),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001110100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46698),
    .in1(net_46699),
    .in2(net_46700_cascademuxed),
    .in3(net_46701),
    .lcout(net_42768),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46704),
    .in1(net_46705),
    .in2(net_46706_cascademuxed),
    .in3(net_46707),
    .lcout(net_42769),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46712_cascademuxed),
    .in3(gnd),
    .lcout(net_42770),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46837),
    .clk(net_46838),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46794),
    .lcout(net_42886),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46798),
    .in2(gnd),
    .in3(net_46800),
    .lcout(net_42887),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46805_cascademuxed),
    .in3(gnd),
    .lcout(net_42888),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46812),
    .lcout(net_42889),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46837),
    .clk(net_46838),
    .in0(net_46815),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42890),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011111110111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46821),
    .in1(net_46822),
    .in2(net_46823_cascademuxed),
    .in3(net_46824),
    .lcout(net_42891),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46837),
    .clk(net_46838),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46829_cascademuxed),
    .in3(gnd),
    .lcout(net_42892),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46833),
    .in1(net_46834),
    .in2(net_46835_cascademuxed),
    .in3(net_46836),
    .lcout(net_42893),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46960),
    .clk(net_46961),
    .in0(gnd),
    .in1(net_46927),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43011),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46932),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43012),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46960),
    .clk(net_46961),
    .in0(gnd),
    .in1(gnd),
    .in2(net_46940_cascademuxed),
    .in3(gnd),
    .lcout(net_43013),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46960),
    .clk(net_46961),
    .in0(gnd),
    .in1(net_46951),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43015),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_11_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47083),
    .clk(net_47084),
    .in0(gnd),
    .in1(gnd),
    .in2(net_47069_cascademuxed),
    .in3(gnd),
    .lcout(net_43137),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_11_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_47207),
    .in0(net_47166),
    .in1(gnd),
    .in2(net_47168_cascademuxed),
    .in3(gnd),
    .lcout(net_43256),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111101110111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_47289),
    .in1(net_47290),
    .in2(net_47291_cascademuxed),
    .in3(net_47292),
    .lcout(net_43379),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010110111111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_47295),
    .in1(net_47296),
    .in2(net_47297_cascademuxed),
    .in3(net_47298),
    .lcout(net_43380),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47329),
    .clk(net_47330),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_47304),
    .lcout(net_43381),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47329),
    .clk(net_47330),
    .in0(gnd),
    .in1(net_47308),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43382),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_11_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47329),
    .clk(net_47330),
    .in0(gnd),
    .in1(net_47314),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43383),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010110111111),
    .SEQ_MODE(4'b0000)
  ) lc40_11_19_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_47418),
    .in1(net_47419),
    .in2(net_47420_cascademuxed),
    .in3(net_47421),
    .lcout(net_43503),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47452),
    .clk(net_47453),
    .in0(net_47424),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43504),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47452),
    .clk(net_47453),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_47445),
    .lcout(net_43507),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47575),
    .clk(net_47576),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_47538),
    .lcout(net_43625),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_20_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47575),
    .clk(net_47576),
    .in0(gnd),
    .in1(gnd),
    .in2(net_47543_cascademuxed),
    .in3(gnd),
    .lcout(net_43626),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_11_20_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47575),
    .clk(net_47576),
    .in0(net_47565),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_43630),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_23_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_47944),
    .clk(net_47945),
    .in0(gnd),
    .in1(gnd),
    .in2(net_47936_cascademuxed),
    .in3(gnd),
    .lcout(net_43999),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_29_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_48668_cascademuxed),
    .in3(net_48669),
    .lcout(net_44736),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101101110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_30_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_48765),
    .in1(net_48766),
    .in2(net_48767_cascademuxed),
    .in3(net_48768),
    .lcout(net_44855),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010001001100),
    .SEQ_MODE(4'b0000)
  ) lc40_11_30_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_48777),
    .in1(net_48778),
    .in2(net_48779_cascademuxed),
    .in3(net_48780),
    .lcout(net_44857),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111001011010000),
    .SEQ_MODE(4'b1000)
  ) lc40_11_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_45976),
    .clk(net_45977),
    .in0(net_45930),
    .in1(net_45931),
    .in2(net_45932_cascademuxed),
    .in3(net_45933),
    .lcout(net_42025),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_7_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_45943),
    .in2(gnd),
    .in3(net_45945),
    .lcout(net_42027),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_45972),
    .in1(gnd),
    .in2(net_45974_cascademuxed),
    .in3(gnd),
    .lcout(net_42032),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_8_0 (
    .carryin(t138),
    .carryout(t140),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46054),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_8_1 (
    .carryin(t140),
    .carryout(net_46058),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46060),
    .in2(net_46061_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_8_2 (
    .carryin(net_46058),
    .carryout(net_46064),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46066),
    .in2(net_46067_cascademuxed),
    .in3(net_46068),
    .lcout(net_42150),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_8_3 (
    .carryin(net_46064),
    .carryout(net_46070),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46072),
    .in2(net_46073_cascademuxed),
    .in3(net_46074),
    .lcout(net_42151),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_8_4 (
    .carryin(net_46070),
    .carryout(net_46076),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46078),
    .in2(net_46079_cascademuxed),
    .in3(net_46080),
    .lcout(net_42152),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_8_5 (
    .carryin(net_46076),
    .carryout(net_46082),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46084),
    .in2(net_46085_cascademuxed),
    .in3(net_46086),
    .lcout(net_42153),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_8_6 (
    .carryin(net_46082),
    .carryout(net_46088),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46090),
    .in2(net_46091_cascademuxed),
    .in3(net_46092),
    .lcout(net_42154),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_11_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46095),
    .in1(gnd),
    .in2(net_46097_cascademuxed),
    .in3(net_46098),
    .lcout(net_42155),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46179),
    .lcout(net_42271),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_46183),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_42272),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_11_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_46197),
    .lcout(net_42274),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010011100110011),
    .SEQ_MODE(4'b1000)
  ) lc40_11_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46222),
    .clk(net_46223),
    .in0(net_46200),
    .in1(net_46201),
    .in2(net_46202_cascademuxed),
    .in3(net_46203),
    .lcout(net_42275),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001101010011),
    .SEQ_MODE(4'b1000)
  ) lc40_11_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46222),
    .clk(net_46223),
    .in0(net_46206),
    .in1(net_46207),
    .in2(net_46208_cascademuxed),
    .in3(net_46209),
    .lcout(net_42276),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101001101010101),
    .SEQ_MODE(4'b1000)
  ) lc40_11_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_46222),
    .clk(net_46223),
    .in0(net_46212),
    .in1(net_46213),
    .in2(net_46214_cascademuxed),
    .in3(net_46215),
    .lcout(net_42277),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_11_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_46218),
    .in1(net_46219),
    .in2(net_46220_cascademuxed),
    .in3(net_46221),
    .lcout(net_42278),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50299),
    .clk(net_50300),
    .in0(net_50253),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46348),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50259),
    .in1(net_50260),
    .in2(net_50261_cascademuxed),
    .in3(net_50262),
    .lcout(net_46349),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50265),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46350),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010011101110111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50271),
    .in1(net_50272),
    .in2(net_50273_cascademuxed),
    .in3(net_50274),
    .lcout(net_46351),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_50284),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46353),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50299),
    .clk(net_50300),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50292),
    .lcout(net_46354),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_12_0 (
    .carryin(t219),
    .carryout(net_50375),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_50377),
    .in2(net_50378_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_1 (
    .carryin(net_50375),
    .carryout(net_50381),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(net_50383),
    .in2(net_50384_cascademuxed),
    .in3(net_50385),
    .lcout(net_46472),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_2 (
    .carryin(net_50381),
    .carryout(net_50387),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(net_50389),
    .in2(net_50390_cascademuxed),
    .in3(net_50391),
    .lcout(net_46473),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_3 (
    .carryin(net_50387),
    .carryout(net_50393),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(net_50395),
    .in2(net_50396_cascademuxed),
    .in3(net_50397),
    .lcout(net_46474),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_4 (
    .carryin(net_50393),
    .carryout(net_50399),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(net_50401),
    .in2(net_50402_cascademuxed),
    .in3(net_50403),
    .lcout(net_46475),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_5 (
    .carryin(net_50399),
    .carryout(net_50405),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(net_50407),
    .in2(net_50408_cascademuxed),
    .in3(net_50409),
    .lcout(net_46476),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_6 (
    .carryin(net_50405),
    .carryout(net_50411),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(net_50413),
    .in2(net_50414_cascademuxed),
    .in3(net_50415),
    .lcout(net_46477),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_12_7 (
    .carryin(net_50411),
    .carryout(net_50417),
    .ce(net_50422),
    .clk(net_50423),
    .in0(gnd),
    .in1(net_50419),
    .in2(net_50420_cascademuxed),
    .in3(net_50421),
    .lcout(net_46478),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_0 (
    .carryin(net_50461),
    .carryout(net_50498),
    .ce(net_50545),
    .clk(net_50546),
    .in0(gnd),
    .in1(net_50500),
    .in2(net_50501_cascademuxed),
    .in3(net_50502),
    .lcout(net_46594),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_1 (
    .carryin(net_50498),
    .carryout(net_50504),
    .ce(net_50545),
    .clk(net_50546),
    .in0(gnd),
    .in1(net_50506),
    .in2(net_50507_cascademuxed),
    .in3(net_50508),
    .lcout(net_46595),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_2 (
    .carryin(net_50504),
    .carryout(net_50510),
    .ce(net_50545),
    .clk(net_50546),
    .in0(gnd),
    .in1(net_50512),
    .in2(net_50513_cascademuxed),
    .in3(net_50514),
    .lcout(net_46596),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_3 (
    .carryin(net_50510),
    .carryout(net_50516),
    .ce(net_50545),
    .clk(net_50546),
    .in0(gnd),
    .in1(net_50518),
    .in2(net_50519_cascademuxed),
    .in3(net_50520),
    .lcout(net_46597),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_4 (
    .carryin(net_50516),
    .carryout(net_50522),
    .ce(net_50545),
    .clk(net_50546),
    .in0(gnd),
    .in1(net_50524),
    .in2(net_50525_cascademuxed),
    .in3(net_50526),
    .lcout(net_46598),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_5 (
    .carryin(net_50522),
    .carryout(net_50528),
    .ce(net_50545),
    .clk(net_50546),
    .in0(gnd),
    .in1(net_50530),
    .in2(net_50531_cascademuxed),
    .in3(net_50532),
    .lcout(net_46599),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_6 (
    .carryin(net_50528),
    .carryout(net_50534),
    .ce(net_50545),
    .clk(net_50546),
    .in0(gnd),
    .in1(net_50536),
    .in2(net_50537_cascademuxed),
    .in3(net_50538),
    .lcout(net_46600),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50545),
    .clk(net_50546),
    .in0(gnd),
    .in1(net_50542),
    .in2(net_50543_cascademuxed),
    .in3(net_50544),
    .lcout(net_46601),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_12_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50668),
    .clk(net_50669),
    .in0(net_50622),
    .in1(net_50623),
    .in2(net_50624_cascademuxed),
    .in3(gnd),
    .lcout(net_46717),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50631),
    .lcout(net_46718),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001101011111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50634),
    .in1(net_50635),
    .in2(net_50636_cascademuxed),
    .in3(net_50637),
    .lcout(net_46719),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50640),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46720),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50649),
    .lcout(net_46721),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50654_cascademuxed),
    .in3(gnd),
    .lcout(net_46722),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001101101011111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50664),
    .in1(net_50665),
    .in2(net_50666_cascademuxed),
    .in3(net_50667),
    .lcout(net_46724),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50791),
    .clk(net_50792),
    .in0(net_50745),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46840),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_50752),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46841),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011111110111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50757),
    .in1(net_50758),
    .in2(net_50759_cascademuxed),
    .in3(net_50760),
    .lcout(net_46842),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50763),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46843),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101001101011111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50769),
    .in1(net_50770),
    .in2(net_50771_cascademuxed),
    .in3(net_50772),
    .lcout(net_46844),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100011101110111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50775),
    .in1(net_50776),
    .in2(net_50777_cascademuxed),
    .in3(net_50778),
    .lcout(net_46845),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50791),
    .clk(net_50792),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50789_cascademuxed),
    .in3(gnd),
    .lcout(net_46847),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50876_cascademuxed),
    .in3(gnd),
    .lcout(net_46964),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50914),
    .clk(net_50915),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_50883),
    .lcout(net_46965),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_50914),
    .clk(net_50915),
    .in0(gnd),
    .in1(net_50893),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46967),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_50898),
    .in1(net_50899),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_46968),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_50905),
    .in2(net_50906_cascademuxed),
    .in3(gnd),
    .lcout(net_46969),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50993_cascademuxed),
    .in3(gnd),
    .lcout(net_47086),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51037),
    .clk(net_51038),
    .in0(gnd),
    .in1(gnd),
    .in2(net_50999_cascademuxed),
    .in3(gnd),
    .lcout(net_47087),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_51012),
    .lcout(net_47089),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51037),
    .clk(net_51038),
    .in0(gnd),
    .in1(net_51022),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47091),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_51027),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47092),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110001111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_51114),
    .in1(net_51115),
    .in2(net_51116_cascademuxed),
    .in3(net_51117),
    .lcout(net_47209),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001101101011111),
    .SEQ_MODE(4'b0000)
  ) lc40_12_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_51126),
    .in1(net_51127),
    .in2(net_51128_cascademuxed),
    .in3(net_51129),
    .lcout(net_47211),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_12_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51160),
    .clk(net_51161),
    .in0(net_51144),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47214),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51160),
    .clk(net_51161),
    .in0(gnd),
    .in1(net_51157),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47216),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110110011),
    .SEQ_MODE(4'b0000)
  ) lc40_12_19_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_51249),
    .in1(net_51250),
    .in2(net_51251_cascademuxed),
    .in3(net_51252),
    .lcout(net_47334),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51283),
    .clk(net_51284),
    .in0(gnd),
    .in1(net_51256),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47335),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_19_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_51261),
    .in1(gnd),
    .in2(net_51263_cascademuxed),
    .in3(gnd),
    .lcout(net_47336),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51283),
    .clk(net_51284),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_51276),
    .lcout(net_47338),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_51280),
    .in2(gnd),
    .in3(net_51282),
    .lcout(net_47339),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51406),
    .clk(net_51407),
    .in0(gnd),
    .in1(net_51367),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47456),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_21_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_51484),
    .in2(net_51485_cascademuxed),
    .in3(gnd),
    .lcout(net_47578),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_21_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_51529),
    .clk(net_51530),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_51498),
    .lcout(net_47580),
    .ltout(),
    .sr(net_51531)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_21_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_51508),
    .in2(gnd),
    .in3(net_51510),
    .lcout(net_47582),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_21_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_51521_cascademuxed),
    .in3(net_51522),
    .lcout(net_47584),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010001010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_12_21_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_51525),
    .in1(net_51526),
    .in2(net_51527_cascademuxed),
    .in3(net_51528),
    .lcout(net_47585),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_23_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_51776),
    .in0(gnd),
    .in1(net_51730),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_47824),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_26_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_27_0 (
    .carryin(t245),
    .carryout(t247),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_52223_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_27_1 (
    .carryin(t247),
    .carryout(net_52226),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_52229_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_12_27_2 (
    .carryin(net_52226),
    .carryout(net_52232),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_52234),
    .in2(gnd),
    .in3(net_52236),
    .lcout(net_48318),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_12_27_3 (
    .carryin(net_52232),
    .carryout(net_52238),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_52241_cascademuxed),
    .in3(net_52242),
    .lcout(net_48319),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_12_27_4 (
    .carryin(net_52238),
    .carryout(net_52244),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_52246),
    .in2(gnd),
    .in3(net_52248),
    .lcout(net_48320),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_12_27_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_52252),
    .in2(gnd),
    .in3(net_52254),
    .lcout(net_48321),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_27_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_52267),
    .clk(net_52268),
    .in0(net_52257),
    .in1(net_52258),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_48322),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_27_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_52267),
    .clk(net_52268),
    .in0(gnd),
    .in1(net_52264),
    .in2(gnd),
    .in3(net_52266),
    .lcout(net_48323),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_12_28_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_52390),
    .clk(net_52391),
    .in0(gnd),
    .in1(gnd),
    .in2(net_52352_cascademuxed),
    .in3(net_52353),
    .lcout(net_48440),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_12_28_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_52356),
    .in1(gnd),
    .in2(net_52358_cascademuxed),
    .in3(gnd),
    .lcout(net_48441),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_12_30_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_48691),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_12_8_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_49892_cascademuxed),
    .in3(gnd),
    .lcout(net_45980),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_12_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_49930),
    .clk(net_49931),
    .in0(gnd),
    .in1(net_49915),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_45984),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000010),
    .SEQ_MODE(4'b0000)
  ) lc40_12_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_49920),
    .in1(gnd),
    .in2(net_49922_cascademuxed),
    .in3(net_49923),
    .lcout(net_45985),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54090),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50180),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54130),
    .clk(net_54131),
    .in0(net_54120),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50185),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011111110111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54207),
    .in1(net_54208),
    .in2(net_54209_cascademuxed),
    .in3(net_54210),
    .lcout(net_50302),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_54214),
    .in2(net_54215_cascademuxed),
    .in3(gnd),
    .lcout(net_50303),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010110111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54219),
    .in1(net_54220),
    .in2(net_54221_cascademuxed),
    .in3(net_54222),
    .lcout(net_50304),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54225),
    .in1(net_54226),
    .in2(net_54227_cascademuxed),
    .in3(net_54228),
    .lcout(net_50305),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54234),
    .lcout(net_50306),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54253),
    .clk(net_54254),
    .in0(gnd),
    .in1(net_54238),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50307),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011111110111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54243),
    .in1(net_54244),
    .in2(net_54245_cascademuxed),
    .in3(net_54246),
    .lcout(net_50308),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54252),
    .lcout(net_50309),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111111001111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54330),
    .in1(net_54331),
    .in2(net_54332_cascademuxed),
    .in3(net_54333),
    .lcout(net_50425),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54338_cascademuxed),
    .in3(gnd),
    .lcout(net_50426),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001111011111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54342),
    .in1(net_54343),
    .in2(net_54344_cascademuxed),
    .in3(net_54345),
    .lcout(net_50427),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54348),
    .in1(net_54349),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50428),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54376),
    .clk(net_54377),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54356_cascademuxed),
    .in3(gnd),
    .lcout(net_50429),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54376),
    .clk(net_54377),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54363),
    .lcout(net_50430),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54376),
    .clk(net_54377),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54369),
    .lcout(net_50431),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54372),
    .in1(net_54373),
    .in2(net_54374_cascademuxed),
    .in3(net_54375),
    .lcout(net_50432),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001110100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54453),
    .in1(net_54454),
    .in2(net_54455_cascademuxed),
    .in3(net_54456),
    .lcout(net_50548),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54459),
    .in1(gnd),
    .in2(net_54461_cascademuxed),
    .in3(gnd),
    .lcout(net_50549),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54467_cascademuxed),
    .in3(gnd),
    .lcout(net_50550),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010110111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54471),
    .in1(net_54472),
    .in2(net_54473_cascademuxed),
    .in3(net_54474),
    .lcout(net_50551),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_54478),
    .in2(gnd),
    .in3(net_54480),
    .lcout(net_50552),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54499),
    .clk(net_54500),
    .in0(net_54483),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50553),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54489),
    .in1(net_54490),
    .in2(net_54491_cascademuxed),
    .in3(net_54492),
    .lcout(net_50554),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54499),
    .clk(net_54500),
    .in0(gnd),
    .in1(net_54496),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50555),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110101011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54576),
    .in1(net_54577),
    .in2(net_54578_cascademuxed),
    .in3(net_54579),
    .lcout(net_50671),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54622),
    .clk(net_54623),
    .in0(net_54582),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50672),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54622),
    .clk(net_54623),
    .in0(gnd),
    .in1(net_54589),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_50673),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_54595),
    .in2(net_54596_cascademuxed),
    .in3(gnd),
    .lcout(net_50674),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54603),
    .lcout(net_50675),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_54609),
    .lcout(net_50676),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_54614_cascademuxed),
    .in3(gnd),
    .lcout(net_50677),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110111011101),
    .SEQ_MODE(4'b0000)
  ) lc40_13_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_54618),
    .in1(net_54619),
    .in2(net_54620_cascademuxed),
    .in3(net_54621),
    .lcout(net_50678),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_16_0 (
    .carryin(t285),
    .carryout(net_54698),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_54700),
    .in2(net_54701_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_1 (
    .carryin(net_54698),
    .carryout(net_54704),
    .ce(net_54745),
    .clk(net_54746),
    .in0(gnd),
    .in1(net_54706),
    .in2(net_54707_cascademuxed),
    .in3(net_54708),
    .lcout(net_50795),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_2 (
    .carryin(net_54704),
    .carryout(net_54710),
    .ce(net_54745),
    .clk(net_54746),
    .in0(gnd),
    .in1(net_54712),
    .in2(net_54713_cascademuxed),
    .in3(net_54714),
    .lcout(net_50796),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_3 (
    .carryin(net_54710),
    .carryout(net_54716),
    .ce(net_54745),
    .clk(net_54746),
    .in0(gnd),
    .in1(net_54718),
    .in2(net_54719_cascademuxed),
    .in3(net_54720),
    .lcout(net_50797),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_4 (
    .carryin(net_54716),
    .carryout(net_54722),
    .ce(net_54745),
    .clk(net_54746),
    .in0(gnd),
    .in1(net_54724),
    .in2(net_54725_cascademuxed),
    .in3(net_54726),
    .lcout(net_50798),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_5 (
    .carryin(net_54722),
    .carryout(net_54728),
    .ce(net_54745),
    .clk(net_54746),
    .in0(gnd),
    .in1(net_54730),
    .in2(net_54731_cascademuxed),
    .in3(net_54732),
    .lcout(net_50799),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_6 (
    .carryin(net_54728),
    .carryout(net_54734),
    .ce(net_54745),
    .clk(net_54746),
    .in0(gnd),
    .in1(net_54736),
    .in2(net_54737_cascademuxed),
    .in3(net_54738),
    .lcout(net_50800),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_16_7 (
    .carryin(net_54734),
    .carryout(net_54740),
    .ce(net_54745),
    .clk(net_54746),
    .in0(gnd),
    .in1(net_54742),
    .in2(net_54743_cascademuxed),
    .in3(net_54744),
    .lcout(net_50801),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_0 (
    .carryin(net_54784),
    .carryout(net_54821),
    .ce(net_54868),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54823),
    .in2(net_54824_cascademuxed),
    .in3(net_54825),
    .lcout(net_50917),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_1 (
    .carryin(net_54821),
    .carryout(net_54827),
    .ce(net_54868),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54829),
    .in2(net_54830_cascademuxed),
    .in3(net_54831),
    .lcout(net_50918),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_2 (
    .carryin(net_54827),
    .carryout(net_54833),
    .ce(net_54868),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54835),
    .in2(net_54836_cascademuxed),
    .in3(net_54837),
    .lcout(net_50919),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_3 (
    .carryin(net_54833),
    .carryout(net_54839),
    .ce(net_54868),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54841),
    .in2(net_54842_cascademuxed),
    .in3(net_54843),
    .lcout(net_50920),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_4 (
    .carryin(net_54839),
    .carryout(net_54845),
    .ce(net_54868),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54847),
    .in2(net_54848_cascademuxed),
    .in3(net_54849),
    .lcout(net_50921),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_5 (
    .carryin(net_54845),
    .carryout(net_54851),
    .ce(net_54868),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54853),
    .in2(net_54854_cascademuxed),
    .in3(net_54855),
    .lcout(net_50922),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_6 (
    .carryin(net_54851),
    .carryout(net_54857),
    .ce(net_54868),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54859),
    .in2(net_54860_cascademuxed),
    .in3(net_54861),
    .lcout(net_50923),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_13_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54868),
    .clk(net_54869),
    .in0(gnd),
    .in1(net_54865),
    .in2(net_54866_cascademuxed),
    .in3(net_54867),
    .lcout(net_50924),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(gnd),
    .in1(net_54964),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_51043),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(gnd),
    .in1(net_54970),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_51044),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_13_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_54991),
    .clk(net_54992),
    .in0(gnd),
    .in1(net_54976),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_51045),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110111110101),
    .SEQ_MODE(4'b0000)
  ) lc40_13_19_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_55074),
    .in1(net_55075),
    .in2(net_55076_cascademuxed),
    .in3(net_55077),
    .lcout(net_51164),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_19_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55114),
    .clk(net_55115),
    .in0(gnd),
    .in1(gnd),
    .in2(net_55082_cascademuxed),
    .in3(gnd),
    .lcout(net_51165),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111100011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_19_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_55092),
    .in1(net_55093),
    .in2(net_55094_cascademuxed),
    .in3(net_55095),
    .lcout(net_51167),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001111011111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_55104),
    .in1(net_55105),
    .in2(net_55106_cascademuxed),
    .in3(net_55107),
    .lcout(net_51169),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55114),
    .clk(net_55115),
    .in0(gnd),
    .in1(gnd),
    .in2(net_55112_cascademuxed),
    .in3(gnd),
    .lcout(net_51170),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_20_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55237),
    .clk(net_55238),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_55194),
    .lcout(net_51286),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55237),
    .clk(net_55238),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_55200),
    .lcout(net_51287),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_20_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55237),
    .clk(net_55238),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_55212),
    .lcout(net_51289),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_20_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55237),
    .clk(net_55238),
    .in0(gnd),
    .in1(gnd),
    .in2(net_55217_cascademuxed),
    .in3(gnd),
    .lcout(net_51290),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_20_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55237),
    .clk(net_55238),
    .in0(gnd),
    .in1(gnd),
    .in2(net_55223_cascademuxed),
    .in3(gnd),
    .lcout(net_51291),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010110111111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_20_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_55227),
    .in1(net_55228),
    .in2(net_55229_cascademuxed),
    .in3(net_55230),
    .lcout(net_51292),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001101011111),
    .SEQ_MODE(4'b0000)
  ) lc40_13_20_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_55233),
    .in1(net_55234),
    .in2(net_55235_cascademuxed),
    .in3(net_55236),
    .lcout(net_51293),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_21_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_55351),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_51415),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_22_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55483),
    .clk(net_55484),
    .in0(net_55443),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_51533),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000001100),
    .SEQ_MODE(4'b0000)
  ) lc40_13_22_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_55455),
    .in1(net_55456),
    .in2(net_55457_cascademuxed),
    .in3(net_55458),
    .lcout(net_51535),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_22_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_55483),
    .clk(net_55484),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_55470),
    .lcout(net_51537),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_22_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_55479),
    .in1(net_55480),
    .in2(net_55481_cascademuxed),
    .in3(net_55482),
    .lcout(net_51539),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_27_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56064),
    .in1(net_56065),
    .in2(net_56066_cascademuxed),
    .in3(net_56067),
    .lcout(net_52149),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_27_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56098),
    .clk(net_56099),
    .in0(net_56076),
    .in1(gnd),
    .in2(gnd),
    .in3(net_56079),
    .lcout(net_52151),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_27_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56098),
    .clk(net_56099),
    .in0(net_56082),
    .in1(gnd),
    .in2(net_56084_cascademuxed),
    .in3(net_56085),
    .lcout(net_52152),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_27_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56088),
    .in1(net_56089),
    .in2(net_56090_cascademuxed),
    .in3(net_56091),
    .lcout(net_52153),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_27_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56098),
    .clk(net_56099),
    .in0(net_56094),
    .in1(net_56095),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_52154),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53146),
    .clk(net_53147),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_53109),
    .lcout(net_49196),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53142),
    .in1(net_53143),
    .in2(net_53144_cascademuxed),
    .in3(net_53145),
    .lcout(net_49202),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_4_0 (
    .carryin(t251),
    .carryout(t253),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53225_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_4_1 (
    .carryin(t253),
    .carryout(net_53228),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53231_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_4_2 (
    .carryin(net_53228),
    .carryout(net_53234),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53237_cascademuxed),
    .in3(net_53238),
    .lcout(net_49320),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_4_3 (
    .carryin(net_53234),
    .carryout(net_53240),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_53242),
    .in2(gnd),
    .in3(net_53244),
    .lcout(net_49321),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_4_4 (
    .carryin(net_53240),
    .carryout(net_53246),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_53248),
    .in2(gnd),
    .in3(net_53250),
    .lcout(net_49322),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53255_cascademuxed),
    .in3(net_53256),
    .lcout(net_49323),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_4_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53269),
    .clk(net_53270),
    .in0(net_53259),
    .in1(net_53260),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_49324),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53269),
    .clk(net_53270),
    .in0(net_53265),
    .in1(gnd),
    .in2(net_53267_cascademuxed),
    .in3(gnd),
    .lcout(net_49325),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_0 (
    .carryin(t254),
    .carryout(t256),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_53716),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_1 (
    .carryin(t256),
    .carryout(net_53720),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_53722),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_2 (
    .carryin(net_53720),
    .carryout(net_53726),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_53728),
    .in2(gnd),
    .in3(net_53730),
    .lcout(net_49812),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_3 (
    .carryin(net_53726),
    .carryout(net_53732),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53735_cascademuxed),
    .in3(net_53736),
    .lcout(net_49813),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_4 (
    .carryin(net_53732),
    .carryout(net_53738),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53741_cascademuxed),
    .in3(net_53742),
    .lcout(net_49814),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_5 (
    .carryin(net_53738),
    .carryout(net_53744),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53747_cascademuxed),
    .in3(net_53748),
    .lcout(net_49815),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_6 (
    .carryin(net_53744),
    .carryout(net_53750),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53753_cascademuxed),
    .in3(net_53754),
    .lcout(net_49816),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_13_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_53759_cascademuxed),
    .in3(net_53760),
    .lcout(net_49817),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011100010101010),
    .SEQ_MODE(4'b1000)
  ) lc40_13_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53884),
    .clk(net_53885),
    .in0(net_53838),
    .in1(net_53839),
    .in2(net_53840_cascademuxed),
    .in3(net_53841),
    .lcout(net_49933),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111101000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53884),
    .clk(net_53885),
    .in0(net_53844),
    .in1(net_53845),
    .in2(net_53846_cascademuxed),
    .in3(net_53847),
    .lcout(net_49934),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_13_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_53850),
    .in1(net_53851),
    .in2(net_53852_cascademuxed),
    .in3(net_53853),
    .lcout(net_49935),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111101000000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53884),
    .clk(net_53885),
    .in0(net_53868),
    .in1(net_53869),
    .in2(net_53870_cascademuxed),
    .in3(net_53871),
    .lcout(net_49938),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110001011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_13_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_53884),
    .clk(net_53885),
    .in0(net_53874),
    .in1(net_53875),
    .in2(net_53876_cascademuxed),
    .in3(net_53877),
    .lcout(net_49939),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57833),
    .in1(net_57834),
    .in2(net_57835_cascademuxed),
    .in3(net_57836),
    .lcout(net_53894),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57915),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54010),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57960),
    .clk(net_57961),
    .in0(net_57920),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54011),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110111011101),
    .SEQ_MODE(4'b0000)
  ) lc40_14_11_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57926),
    .in1(net_57927),
    .in2(net_57928_cascademuxed),
    .in3(net_57929),
    .lcout(net_54012),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_11_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57960),
    .clk(net_57961),
    .in0(gnd),
    .in1(net_57933),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54013),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001101011111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57938),
    .in1(net_57939),
    .in2(net_57940_cascademuxed),
    .in3(net_57941),
    .lcout(net_54014),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57944),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54015),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_11_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57952_cascademuxed),
    .in3(gnd),
    .lcout(net_54016),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57960),
    .clk(net_57961),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_57959),
    .lcout(net_54017),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58037),
    .in1(net_58038),
    .in2(net_58039_cascademuxed),
    .in3(net_58040),
    .lcout(net_54133),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58083),
    .clk(net_58084),
    .in0(net_58043),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54134),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001101011111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58049),
    .in1(net_58050),
    .in2(net_58051_cascademuxed),
    .in3(net_58052),
    .lcout(net_54135),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58055),
    .in1(net_58056),
    .in2(net_58057_cascademuxed),
    .in3(net_58058),
    .lcout(net_54136),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58064),
    .lcout(net_54137),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58067),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54138),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58083),
    .clk(net_58084),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58076),
    .lcout(net_54139),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101110111011),
    .SEQ_MODE(4'b0000)
  ) lc40_14_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58079),
    .in1(net_58080),
    .in2(net_58081_cascademuxed),
    .in3(net_58082),
    .lcout(net_54140),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58160),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54256),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111111001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58166),
    .in1(net_58167),
    .in2(net_58168_cascademuxed),
    .in3(net_58169),
    .lcout(net_54257),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001111011111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58172),
    .in1(net_58173),
    .in2(net_58174_cascademuxed),
    .in3(net_58175),
    .lcout(net_54258),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110101011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58178),
    .in1(net_58179),
    .in2(net_58180_cascademuxed),
    .in3(net_58181),
    .lcout(net_54259),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58184),
    .in1(net_58185),
    .in2(net_58186_cascademuxed),
    .in3(net_58187),
    .lcout(net_54260),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110111011101),
    .SEQ_MODE(4'b0000)
  ) lc40_14_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58190),
    .in1(net_58191),
    .in2(net_58192_cascademuxed),
    .in3(net_58193),
    .lcout(net_54261),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101111110011),
    .SEQ_MODE(4'b0000)
  ) lc40_14_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58196),
    .in1(net_58197),
    .in2(net_58198_cascademuxed),
    .in3(net_58199),
    .lcout(net_54262),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58206),
    .clk(net_58207),
    .in0(gnd),
    .in1(net_58203),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54263),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111111001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58283),
    .in1(net_58284),
    .in2(net_58285_cascademuxed),
    .in3(net_58286),
    .lcout(net_54379),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58290),
    .in2(net_58291_cascademuxed),
    .in3(gnd),
    .lcout(net_54380),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110111011101),
    .SEQ_MODE(4'b0000)
  ) lc40_14_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58295),
    .in1(net_58296),
    .in2(net_58297_cascademuxed),
    .in3(net_58298),
    .lcout(net_54381),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58302),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54382),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58309_cascademuxed),
    .in3(net_58310),
    .lcout(net_54383),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58329),
    .clk(net_58330),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58315_cascademuxed),
    .in3(gnd),
    .lcout(net_54384),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58329),
    .clk(net_58330),
    .in0(net_58319),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54385),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111111001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58325),
    .in1(net_58326),
    .in2(net_58327_cascademuxed),
    .in3(net_58328),
    .lcout(net_54386),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58452),
    .clk(net_58453),
    .in0(gnd),
    .in1(net_58407),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54502),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58414_cascademuxed),
    .in3(net_58415),
    .lcout(net_54503),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58452),
    .clk(net_58453),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58420_cascademuxed),
    .in3(gnd),
    .lcout(net_54504),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58424),
    .in1(net_58425),
    .in2(net_58426_cascademuxed),
    .in3(net_58427),
    .lcout(net_54505),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58452),
    .clk(net_58453),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58432_cascademuxed),
    .in3(gnd),
    .lcout(net_54506),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58437),
    .in2(net_58438_cascademuxed),
    .in3(gnd),
    .lcout(net_54507),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58452),
    .clk(net_58453),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58445),
    .lcout(net_54508),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58452),
    .clk(net_58453),
    .in0(net_58448),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54509),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_58531_cascademuxed),
    .in3(gnd),
    .lcout(net_54625),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58535),
    .in1(net_58536),
    .in2(net_58537_cascademuxed),
    .in3(net_58538),
    .lcout(net_54626),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58550),
    .lcout(net_54628),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58553),
    .in1(gnd),
    .in2(net_58555_cascademuxed),
    .in3(gnd),
    .lcout(net_54629),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58575),
    .clk(net_58576),
    .in0(net_58559),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54630),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58568),
    .lcout(net_54631),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58571),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54632),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58698),
    .clk(net_58699),
    .in0(net_58658),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54749),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58665),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54750),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58671),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54751),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58682),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58685),
    .lcout(net_54753),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58695),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54755),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58776),
    .in2(gnd),
    .in3(net_58778),
    .lcout(net_54871),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(net_58781),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54872),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58793),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58796),
    .lcout(net_54874),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58799),
    .in1(net_58800),
    .in2(net_58801_cascademuxed),
    .in3(net_58802),
    .lcout(net_54875),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58821),
    .clk(net_58822),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_58808),
    .lcout(net_54876),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110001111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58817),
    .in1(net_58818),
    .in2(net_58819_cascademuxed),
    .in3(net_58820),
    .lcout(net_54878),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_19_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_58944),
    .clk(net_58945),
    .in0(gnd),
    .in1(net_58899),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_54994),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_19_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_58904),
    .in1(net_58905),
    .in2(net_58906_cascademuxed),
    .in3(net_58907),
    .lcout(net_54995),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58935),
    .in2(net_58936_cascademuxed),
    .in3(gnd),
    .lcout(net_55000),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_58941),
    .in2(gnd),
    .in3(net_58943),
    .lcout(net_55001),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_20_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_59067),
    .clk(net_59068),
    .in0(gnd),
    .in1(gnd),
    .in2(net_59023_cascademuxed),
    .in3(gnd),
    .lcout(net_55117),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_59027),
    .in1(gnd),
    .in2(net_59029_cascademuxed),
    .in3(gnd),
    .lcout(net_55118),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_20_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_59067),
    .clk(net_59068),
    .in0(gnd),
    .in1(gnd),
    .in2(net_59035_cascademuxed),
    .in3(gnd),
    .lcout(net_55119),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_20_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_59067),
    .clk(net_59068),
    .in0(gnd),
    .in1(net_59046),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_55121),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101110111011),
    .SEQ_MODE(4'b0000)
  ) lc40_14_20_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_59051),
    .in1(net_59052),
    .in2(net_59053_cascademuxed),
    .in3(net_59054),
    .lcout(net_55122),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011111110111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_20_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_59063),
    .in1(net_59064),
    .in2(net_59065_cascademuxed),
    .in3(net_59066),
    .lcout(net_55124),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_21_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_59190),
    .clk(net_59191),
    .in0(gnd),
    .in1(net_59187),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_55247),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_26_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_59805),
    .clk(net_59806),
    .in0(gnd),
    .in1(net_59778),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_55858),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b0000)
  ) lc40_14_26_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_59783),
    .in1(gnd),
    .in2(net_59785_cascademuxed),
    .in3(gnd),
    .lcout(net_55859),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010011101000101),
    .SEQ_MODE(4'b1000)
  ) lc40_14_27_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_59928),
    .clk(net_59929),
    .in0(net_59888),
    .in1(net_59889),
    .in2(net_59890_cascademuxed),
    .in3(net_59891),
    .lcout(net_55979),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_27_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_59895),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_55980),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_27_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_59913),
    .in2(net_59914_cascademuxed),
    .in3(net_59915),
    .lcout(net_55983),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b0000)
  ) lc40_14_28_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_60011),
    .in1(gnd),
    .in2(gnd),
    .in3(net_60014),
    .lcout(net_56102),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56819),
    .in1(gnd),
    .in2(net_56821_cascademuxed),
    .in3(gnd),
    .lcout(net_52869),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110010010101),
    .SEQ_MODE(4'b0000)
  ) lc40_14_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56825),
    .in1(net_56826),
    .in2(net_56827_cascademuxed),
    .in3(net_56828),
    .lcout(net_52870),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010001010000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_56838),
    .in2(net_56839_cascademuxed),
    .in3(net_56840),
    .lcout(net_52872),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56843),
    .in1(net_56844),
    .in2(net_56845_cascademuxed),
    .in3(net_56846),
    .lcout(net_52873),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56930),
    .in1(net_56931),
    .in2(net_56932_cascademuxed),
    .in3(net_56933),
    .lcout(net_53026),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_56937),
    .in2(net_56938_cascademuxed),
    .in3(net_56939),
    .lcout(net_53027),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56942),
    .in1(net_56943),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53028),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1001100001011101),
    .SEQ_MODE(4'b1000)
  ) lc40_14_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_56976),
    .clk(net_56977),
    .in0(net_56948),
    .in1(net_56949),
    .in2(net_56950_cascademuxed),
    .in3(net_56951),
    .lcout(net_53029),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_14_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56954),
    .in1(net_56955),
    .in2(net_56956_cascademuxed),
    .in3(net_56957),
    .lcout(net_53030),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111111110010),
    .SEQ_MODE(4'b0000)
  ) lc40_14_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56960),
    .in1(net_56961),
    .in2(net_56962_cascademuxed),
    .in3(net_56963),
    .lcout(net_53031),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110101111111111),
    .SEQ_MODE(4'b0000)
  ) lc40_14_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56966),
    .in1(net_56967),
    .in2(net_56968_cascademuxed),
    .in3(net_56969),
    .lcout(net_53032),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_56972),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_53033),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(net_57053),
    .in1(net_57054),
    .in2(gnd),
    .in3(net_57056),
    .lcout(net_53149),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(net_57059),
    .in1(gnd),
    .in2(net_57061_cascademuxed),
    .in3(gnd),
    .lcout(net_53150),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_4_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57066),
    .in2(gnd),
    .in3(net_57068),
    .lcout(net_53151),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(gnd),
    .in1(net_57078),
    .in2(gnd),
    .in3(net_57080),
    .lcout(net_53153),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57083),
    .in1(gnd),
    .in2(net_57085_cascademuxed),
    .in3(gnd),
    .lcout(net_53154),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57099),
    .clk(net_57100),
    .in0(gnd),
    .in1(gnd),
    .in2(net_57097_cascademuxed),
    .in3(net_57098),
    .lcout(net_53156),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_7_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57428),
    .in1(gnd),
    .in2(net_57430_cascademuxed),
    .in3(gnd),
    .lcout(net_53519),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_14_7_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57468),
    .clk(net_57469),
    .in0(net_57458),
    .in1(net_57459),
    .in2(net_57460_cascademuxed),
    .in3(net_57461),
    .lcout(net_53524),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57464),
    .in1(gnd),
    .in2(net_57466_cascademuxed),
    .in3(gnd),
    .lcout(net_53525),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_14_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57569),
    .in1(net_57570),
    .in2(net_57571_cascademuxed),
    .in3(net_57572),
    .lcout(net_53645),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100001000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57575),
    .in1(net_57576),
    .in2(gnd),
    .in3(net_57578),
    .lcout(net_53646),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111100100000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57591),
    .clk(net_57592),
    .in0(net_57581),
    .in1(net_57582),
    .in2(net_57583_cascademuxed),
    .in3(net_57584),
    .lcout(net_53647),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_14_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_57591),
    .clk(net_57592),
    .in0(net_57587),
    .in1(net_57588),
    .in2(net_57589_cascademuxed),
    .in3(net_57590),
    .lcout(net_53648),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_0 (
    .carryin(t315),
    .carryout(t317),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57669),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_1 (
    .carryin(t317),
    .carryout(net_57673),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57675),
    .in2(net_57676_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_2 (
    .carryin(net_57673),
    .carryout(net_57679),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57681),
    .in2(net_57682_cascademuxed),
    .in3(net_57683),
    .lcout(net_53766),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_3 (
    .carryin(net_57679),
    .carryout(net_57685),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57687),
    .in2(net_57688_cascademuxed),
    .in3(net_57689),
    .lcout(net_53767),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_4 (
    .carryin(net_57685),
    .carryout(net_57691),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57693),
    .in2(net_57694_cascademuxed),
    .in3(net_57695),
    .lcout(net_53768),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_5 (
    .carryin(net_57691),
    .carryout(net_57697),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57699),
    .in2(net_57700_cascademuxed),
    .in3(net_57701),
    .lcout(net_53769),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_6 (
    .carryin(net_57697),
    .carryout(net_57703),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_57705),
    .in2(net_57706_cascademuxed),
    .in3(net_57707),
    .lcout(net_53770),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_14_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_57710),
    .in1(gnd),
    .in2(net_57712_cascademuxed),
    .in3(net_57713),
    .lcout(net_53771),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_10_0 (
    .carryin(t455),
    .carryout(t458),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61623_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_10_1 (
    .carryin(t458),
    .carryout(net_61626),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61629_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_15_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_61634),
    .in2(gnd),
    .in3(net_61636),
    .lcout(net_57719),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b0000)
  ) lc40_15_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_61645),
    .in1(net_61646),
    .in2(net_61647_cascademuxed),
    .in3(net_61648),
    .lcout(net_57721),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100110000001100),
    .SEQ_MODE(4'b0000)
  ) lc40_15_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_61651),
    .in1(net_61652),
    .in2(net_61653_cascademuxed),
    .in3(net_61654),
    .lcout(net_57722),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61667),
    .clk(net_61668),
    .in0(net_61657),
    .in1(net_61658),
    .in2(net_61659_cascademuxed),
    .in3(gnd),
    .lcout(net_57723),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_11_0 (
    .carryin(t399),
    .carryout(net_61743),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_61745),
    .in2(net_61746_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_1 (
    .carryin(net_61743),
    .carryout(net_61749),
    .ce(net_61790),
    .clk(net_61791),
    .in0(gnd),
    .in1(net_61751),
    .in2(net_61752_cascademuxed),
    .in3(net_61753),
    .lcout(net_57841),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_2 (
    .carryin(net_61749),
    .carryout(net_61755),
    .ce(net_61790),
    .clk(net_61791),
    .in0(gnd),
    .in1(net_61757),
    .in2(net_61758_cascademuxed),
    .in3(net_61759),
    .lcout(net_57842),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_3 (
    .carryin(net_61755),
    .carryout(net_61761),
    .ce(net_61790),
    .clk(net_61791),
    .in0(gnd),
    .in1(net_61763),
    .in2(net_61764_cascademuxed),
    .in3(net_61765),
    .lcout(net_57843),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_4 (
    .carryin(net_61761),
    .carryout(net_61767),
    .ce(net_61790),
    .clk(net_61791),
    .in0(gnd),
    .in1(net_61769),
    .in2(net_61770_cascademuxed),
    .in3(net_61771),
    .lcout(net_57844),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_5 (
    .carryin(net_61767),
    .carryout(net_61773),
    .ce(net_61790),
    .clk(net_61791),
    .in0(gnd),
    .in1(net_61775),
    .in2(net_61776_cascademuxed),
    .in3(net_61777),
    .lcout(net_57845),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_6 (
    .carryin(net_61773),
    .carryout(net_61779),
    .ce(net_61790),
    .clk(net_61791),
    .in0(gnd),
    .in1(net_61781),
    .in2(net_61782_cascademuxed),
    .in3(net_61783),
    .lcout(net_57846),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_11_7 (
    .carryin(net_61779),
    .carryout(net_61785),
    .ce(net_61790),
    .clk(net_61791),
    .in0(gnd),
    .in1(net_61787),
    .in2(net_61788_cascademuxed),
    .in3(net_61789),
    .lcout(net_57847),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_0 (
    .carryin(net_61829),
    .carryout(net_61866),
    .ce(net_61913),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61868),
    .in2(net_61869_cascademuxed),
    .in3(net_61870),
    .lcout(net_57963),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_1 (
    .carryin(net_61866),
    .carryout(net_61872),
    .ce(net_61913),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61874),
    .in2(net_61875_cascademuxed),
    .in3(net_61876),
    .lcout(net_57964),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_2 (
    .carryin(net_61872),
    .carryout(net_61878),
    .ce(net_61913),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61880),
    .in2(net_61881_cascademuxed),
    .in3(net_61882),
    .lcout(net_57965),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_3 (
    .carryin(net_61878),
    .carryout(net_61884),
    .ce(net_61913),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61886),
    .in2(net_61887_cascademuxed),
    .in3(net_61888),
    .lcout(net_57966),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_4 (
    .carryin(net_61884),
    .carryout(net_61890),
    .ce(net_61913),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61892),
    .in2(net_61893_cascademuxed),
    .in3(net_61894),
    .lcout(net_57967),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_5 (
    .carryin(net_61890),
    .carryout(net_61896),
    .ce(net_61913),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61898),
    .in2(net_61899_cascademuxed),
    .in3(net_61900),
    .lcout(net_57968),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_6 (
    .carryin(net_61896),
    .carryout(net_61902),
    .ce(net_61913),
    .clk(net_61914),
    .in0(gnd),
    .in1(net_61904),
    .in2(net_61905_cascademuxed),
    .in3(net_61906),
    .lcout(net_57969),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61913),
    .clk(net_61914),
    .in0(net_61909),
    .in1(gnd),
    .in2(net_61911_cascademuxed),
    .in3(net_61912),
    .lcout(net_57970),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111010101),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_61990),
    .in1(net_61991),
    .in2(net_61992_cascademuxed),
    .in3(net_61993),
    .lcout(net_58086),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_61996),
    .in1(net_61997),
    .in2(net_61998_cascademuxed),
    .in3(net_61999),
    .lcout(net_58087),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111111001111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62002),
    .in1(net_62003),
    .in2(net_62004_cascademuxed),
    .in3(net_62005),
    .lcout(net_58088),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62010_cascademuxed),
    .in3(gnd),
    .lcout(net_58089),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62017),
    .lcout(net_58090),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111010101),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62020),
    .in1(net_62021),
    .in2(net_62022_cascademuxed),
    .in3(net_62023),
    .lcout(net_58091),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110111011101),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62026),
    .in1(net_62027),
    .in2(net_62028_cascademuxed),
    .in3(net_62029),
    .lcout(net_58092),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_62033),
    .in2(net_62034_cascademuxed),
    .in3(gnd),
    .lcout(net_58093),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62159),
    .clk(net_62160),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62116),
    .lcout(net_58209),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101110111011),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62119),
    .in1(net_62120),
    .in2(net_62121_cascademuxed),
    .in3(net_62122),
    .lcout(net_58210),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62125),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58211),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_62132),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58212),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101111110011),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62137),
    .in1(net_62138),
    .in2(net_62139_cascademuxed),
    .in3(net_62140),
    .lcout(net_58213),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62159),
    .clk(net_62160),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62145_cascademuxed),
    .in3(gnd),
    .lcout(net_58214),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62149),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58215),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62155),
    .in1(net_62156),
    .in2(net_62157_cascademuxed),
    .in3(net_62158),
    .lcout(net_58216),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62282),
    .clk(net_62283),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62239),
    .lcout(net_58332),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62282),
    .clk(net_62283),
    .in0(gnd),
    .in1(net_62243),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58333),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110101011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62248),
    .in1(net_62249),
    .in2(net_62250_cascademuxed),
    .in3(net_62251),
    .lcout(net_58334),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62256_cascademuxed),
    .in3(gnd),
    .lcout(net_58335),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111100011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62260),
    .in1(net_62261),
    .in2(net_62262_cascademuxed),
    .in3(net_62263),
    .lcout(net_58336),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62266),
    .in1(gnd),
    .in2(net_62268_cascademuxed),
    .in3(gnd),
    .lcout(net_58337),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62275),
    .lcout(net_58338),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62282),
    .clk(net_62283),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62280_cascademuxed),
    .in3(gnd),
    .lcout(net_58339),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_16_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62359),
    .in1(net_62360),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58455),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62377),
    .in1(net_62378),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58458),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62383),
    .in1(net_62384),
    .in2(net_62385_cascademuxed),
    .in3(net_62386),
    .lcout(net_58459),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_16_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62392),
    .lcout(net_58460),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_15_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62405),
    .clk(net_62406),
    .in0(net_62395),
    .in1(net_62396),
    .in2(gnd),
    .in3(net_62398),
    .lcout(net_58461),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_62402),
    .in2(net_62403_cascademuxed),
    .in3(gnd),
    .lcout(net_58462),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62528),
    .clk(net_62529),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62484_cascademuxed),
    .in3(gnd),
    .lcout(net_58578),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62488),
    .in1(net_62489),
    .in2(net_62490_cascademuxed),
    .in3(net_62491),
    .lcout(net_58579),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62528),
    .clk(net_62529),
    .in0(gnd),
    .in1(net_62495),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58580),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62502_cascademuxed),
    .in3(net_62503),
    .lcout(net_58581),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_62513),
    .in2(gnd),
    .in3(net_62515),
    .lcout(net_58583),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_62519),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58584),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62528),
    .clk(net_62529),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62526_cascademuxed),
    .in3(gnd),
    .lcout(net_58585),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101111110011),
    .SEQ_MODE(4'b0000)
  ) lc40_15_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62605),
    .in1(net_62606),
    .in2(net_62607_cascademuxed),
    .in3(net_62608),
    .lcout(net_58701),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62611),
    .in1(net_62612),
    .in2(net_62613_cascademuxed),
    .in3(net_62614),
    .lcout(net_58702),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62651),
    .clk(net_62652),
    .in0(gnd),
    .in1(gnd),
    .in2(net_62619_cascademuxed),
    .in3(gnd),
    .lcout(net_58703),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62651),
    .clk(net_62652),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62632),
    .lcout(net_58705),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111111001111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62641),
    .in1(net_62642),
    .in2(net_62643_cascademuxed),
    .in3(net_62644),
    .lcout(net_58707),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62651),
    .clk(net_62652),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62650),
    .lcout(net_58708),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_19_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62774),
    .clk(net_62775),
    .in0(gnd),
    .in1(net_62729),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58824),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62746),
    .in1(net_62747),
    .in2(net_62748_cascademuxed),
    .in3(gnd),
    .lcout(net_58827),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_19_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62774),
    .clk(net_62775),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_62761),
    .lcout(net_58829),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62764),
    .in1(gnd),
    .in2(net_62766_cascademuxed),
    .in3(gnd),
    .lcout(net_58830),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_20_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_62897),
    .clk(net_62898),
    .in0(net_62851),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_58947),
    .ltout(),
    .sr(net_62899)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_20_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62863),
    .in1(gnd),
    .in2(net_62865_cascademuxed),
    .in3(gnd),
    .lcout(net_58949),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100010101010),
    .SEQ_MODE(4'b0000)
  ) lc40_15_20_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_62887),
    .in1(net_62888),
    .in2(net_62889_cascademuxed),
    .in3(net_62890),
    .lcout(net_58953),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_20_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_62894),
    .in2(net_62895_cascademuxed),
    .in3(gnd),
    .lcout(net_58954),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_21_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63010),
    .in1(net_63011),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_59076),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_22_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63121),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_59197),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_22_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_63143),
    .clk(net_63144),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_63130),
    .lcout(net_59198),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_23_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_63266),
    .clk(net_63267),
    .in0(gnd),
    .in1(gnd),
    .in2(net_63228_cascademuxed),
    .in3(gnd),
    .lcout(net_59317),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000101010),
    .SEQ_MODE(4'b0000)
  ) lc40_15_23_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63250),
    .in1(net_63251),
    .in2(net_63252_cascademuxed),
    .in3(net_63253),
    .lcout(net_59321),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_23_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63262),
    .in1(net_63263),
    .in2(net_63264_cascademuxed),
    .in3(net_63265),
    .lcout(net_59323),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_25_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_63512),
    .clk(net_63513),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_63499),
    .lcout(net_59567),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_27_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_63743),
    .in2(gnd),
    .in3(net_63745),
    .lcout(net_59813),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110111110111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_28_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63835),
    .in1(net_63836),
    .in2(net_63837_cascademuxed),
    .in3(net_63838),
    .lcout(net_59931),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_28_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63841),
    .in1(net_63842),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_59932),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_28_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63859),
    .in1(net_63860),
    .in2(net_63861_cascademuxed),
    .in3(net_63862),
    .lcout(net_59935),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_28_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63865),
    .in1(net_63866),
    .in2(net_63867_cascademuxed),
    .in3(net_63868),
    .lcout(net_59936),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_28_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63877),
    .in1(net_63878),
    .in2(net_63879_cascademuxed),
    .in3(net_63880),
    .lcout(net_59938),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111100010010101),
    .SEQ_MODE(4'b0000)
  ) lc40_15_29_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_63988),
    .in1(net_63989),
    .in2(net_63990_cascademuxed),
    .in3(net_63991),
    .lcout(net_60059),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_29_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64001),
    .in2(net_64002_cascademuxed),
    .in3(net_64003),
    .lcout(net_60061),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010010),
    .SEQ_MODE(4'b1000)
  ) lc40_15_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_60683),
    .clk(net_60684),
    .in0(net_60637),
    .in1(net_60638),
    .in2(net_60639_cascademuxed),
    .in3(gnd),
    .lcout(net_56697),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_60643),
    .in1(net_60644),
    .in2(net_60645_cascademuxed),
    .in3(net_60646),
    .lcout(net_56698),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011011100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_60649),
    .in1(net_60650),
    .in2(net_60651_cascademuxed),
    .in3(net_60652),
    .lcout(net_56699),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001111100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_60655),
    .in1(net_60656),
    .in2(net_60657_cascademuxed),
    .in3(net_60658),
    .lcout(net_56700),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_60673),
    .in1(gnd),
    .in2(gnd),
    .in3(net_60676),
    .lcout(net_56703),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_60767),
    .in2(net_60768_cascademuxed),
    .in3(net_60769),
    .lcout(net_56857),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000111),
    .SEQ_MODE(4'b1000)
  ) lc40_15_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_60806),
    .clk(net_60807),
    .in0(net_60772),
    .in1(net_60773),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_56858),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010100001101),
    .SEQ_MODE(4'b1000)
  ) lc40_15_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_60806),
    .clk(net_60807),
    .in0(net_60778),
    .in1(net_60779),
    .in2(gnd),
    .in3(net_60781),
    .lcout(net_56859),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111010011110111),
    .SEQ_MODE(4'b0000)
  ) lc40_15_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_60784),
    .in1(net_60785),
    .in2(net_60786_cascademuxed),
    .in3(net_60787),
    .lcout(net_56860),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_60791),
    .in2(net_60792_cascademuxed),
    .in3(net_60793),
    .lcout(net_56861),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_60796),
    .in1(net_60797),
    .in2(net_60798_cascademuxed),
    .in3(net_60799),
    .lcout(net_56862),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010000000001100),
    .SEQ_MODE(4'b1000)
  ) lc40_15_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_60806),
    .clk(net_60807),
    .in0(net_60802),
    .in1(net_60803),
    .in2(net_60804_cascademuxed),
    .in3(net_60805),
    .lcout(net_56863),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61175),
    .clk(net_61176),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_61144),
    .lcout(net_57227),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_15_8_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61421),
    .clk(net_61422),
    .in0(gnd),
    .in1(net_61376),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_57471),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_15_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_61498),
    .in1(gnd),
    .in2(gnd),
    .in3(net_61501),
    .lcout(net_57594),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_15_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_61544),
    .clk(net_61545),
    .in0(gnd),
    .in1(gnd),
    .in2(net_61530_cascademuxed),
    .in3(gnd),
    .lcout(net_57599),
    .ltout(),
    .sr(net_61546)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_15_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_61540),
    .in1(gnd),
    .in2(net_61542_cascademuxed),
    .in3(gnd),
    .lcout(net_57601),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_16_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65485),
    .lcout(net_61552),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_16_11_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65576),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61670),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_16_11_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65583_cascademuxed),
    .in3(gnd),
    .lcout(net_61671),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_16_11_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65600),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61674),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65621),
    .clk(net_65622),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65608),
    .lcout(net_61675),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110110011),
    .SEQ_MODE(4'b0000)
  ) lc40_16_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65698),
    .in1(net_65699),
    .in2(net_65700_cascademuxed),
    .in3(net_65701),
    .lcout(net_61793),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111100011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65704),
    .in1(net_65705),
    .in2(net_65706_cascademuxed),
    .in3(net_65707),
    .lcout(net_61794),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65744),
    .clk(net_65745),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65712_cascademuxed),
    .in3(gnd),
    .lcout(net_61795),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_16_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65723),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61797),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65728),
    .in1(net_65729),
    .in2(net_65730_cascademuxed),
    .in3(net_65731),
    .lcout(net_61798),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110110011),
    .SEQ_MODE(4'b0000)
  ) lc40_16_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65734),
    .in1(net_65735),
    .in2(net_65736_cascademuxed),
    .in3(net_65737),
    .lcout(net_61799),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_16_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65868),
    .in0(net_65821),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61916),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111100011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65833),
    .in1(net_65834),
    .in2(net_65835_cascademuxed),
    .in3(net_65836),
    .lcout(net_61918),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_65868),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65842),
    .lcout(net_61919),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_65846),
    .in2(gnd),
    .in3(net_65848),
    .lcout(net_61920),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65952_cascademuxed),
    .in3(net_65953),
    .lcout(net_62040),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65974),
    .in1(gnd),
    .in2(net_65976_cascademuxed),
    .in3(gnd),
    .lcout(net_62044),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65990),
    .clk(net_65991),
    .in0(gnd),
    .in1(net_65987),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62046),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_66068),
    .in2(net_66069_cascademuxed),
    .in3(gnd),
    .lcout(net_62162),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101110111011),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66079),
    .in1(net_66080),
    .in2(net_66081_cascademuxed),
    .in3(net_66082),
    .lcout(net_62164),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66085),
    .in1(gnd),
    .in2(net_66087_cascademuxed),
    .in3(gnd),
    .lcout(net_62165),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66091),
    .in1(gnd),
    .in2(gnd),
    .in3(net_66094),
    .lcout(net_62166),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101110111011),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66097),
    .in1(net_66098),
    .in2(net_66099_cascademuxed),
    .in3(net_66100),
    .lcout(net_62167),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110111110101),
    .SEQ_MODE(4'b0000)
  ) lc40_16_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66103),
    .in1(net_66104),
    .in2(net_66105_cascademuxed),
    .in3(net_66106),
    .lcout(net_62168),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66113),
    .clk(net_66114),
    .in0(gnd),
    .in1(net_66110),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62169),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66196),
    .in1(gnd),
    .in2(net_66198_cascademuxed),
    .in3(gnd),
    .lcout(net_62286),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66236),
    .clk(net_66237),
    .in0(gnd),
    .in1(net_66203),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62287),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66359),
    .clk(net_66360),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66321_cascademuxed),
    .in3(gnd),
    .lcout(net_62409),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66448),
    .in1(net_66449),
    .in2(net_66450_cascademuxed),
    .in3(net_66451),
    .lcout(net_62533),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66482),
    .clk(net_66483),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66456_cascademuxed),
    .in3(gnd),
    .lcout(net_62534),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66460),
    .in1(gnd),
    .in2(gnd),
    .in3(net_66463),
    .lcout(net_62535),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001111011111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_19_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66565),
    .in1(net_66566),
    .in2(net_66567_cascademuxed),
    .in3(net_66568),
    .lcout(net_62655),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_16_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66605),
    .clk(net_66606),
    .in0(net_66577),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62657),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_19_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66605),
    .clk(net_66606),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66585_cascademuxed),
    .in3(gnd),
    .lcout(net_62658),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001110100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_19_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66589),
    .in1(net_66590),
    .in2(net_66591_cascademuxed),
    .in3(net_66592),
    .lcout(net_62659),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_66596),
    .in2(net_66597_cascademuxed),
    .in3(gnd),
    .lcout(net_62660),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_16_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66605),
    .clk(net_66606),
    .in0(net_66601),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62661),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66728),
    .clk(net_66729),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66690_cascademuxed),
    .in3(gnd),
    .lcout(net_62778),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_20_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66728),
    .clk(net_66729),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66696_cascademuxed),
    .in3(gnd),
    .lcout(net_62779),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010100111111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_20_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66700),
    .in1(net_66701),
    .in2(net_66702_cascademuxed),
    .in3(net_66703),
    .lcout(net_62780),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_20_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66728),
    .clk(net_66729),
    .in0(gnd),
    .in1(gnd),
    .in2(net_66708_cascademuxed),
    .in3(gnd),
    .lcout(net_62781),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011111110111),
    .SEQ_MODE(4'b0000)
  ) lc40_16_20_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_66712),
    .in1(net_66713),
    .in2(net_66714_cascademuxed),
    .in3(net_66715),
    .lcout(net_62782),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_16_20_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66728),
    .clk(net_66729),
    .in0(net_66724),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_62784),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_21_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_66851),
    .clk(net_66852),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_66850),
    .lcout(net_62907),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111111011100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_28_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_67712),
    .clk(net_67713),
    .in0(net_67672),
    .in1(net_67673),
    .in2(net_67674_cascademuxed),
    .in3(net_67675),
    .lcout(net_63762),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011110110111100),
    .SEQ_MODE(4'b0000)
  ) lc40_16_28_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_67678),
    .in1(net_67679),
    .in2(net_67680_cascademuxed),
    .in3(net_67681),
    .lcout(net_63763),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010110000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_28_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_67712),
    .clk(net_67713),
    .in0(net_67684),
    .in1(net_67685),
    .in2(net_67686_cascademuxed),
    .in3(net_67687),
    .lcout(net_63764),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_16_28_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_67691),
    .in2(gnd),
    .in3(net_67693),
    .lcout(net_63765),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001101010),
    .SEQ_MODE(4'b1000)
  ) lc40_16_28_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_67712),
    .clk(net_67713),
    .in0(net_67696),
    .in1(net_67697),
    .in2(net_67698_cascademuxed),
    .in3(net_67699),
    .lcout(net_63766),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1011101011101010),
    .SEQ_MODE(4'b1000)
  ) lc40_16_28_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_67712),
    .clk(net_67713),
    .in0(net_67702),
    .in1(net_67703),
    .in2(net_67704_cascademuxed),
    .in3(net_67705),
    .lcout(net_63767),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100100010001000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_28_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_67708),
    .in1(net_67709),
    .in2(net_67710_cascademuxed),
    .in3(net_67711),
    .lcout(net_63768),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110011001011),
    .SEQ_MODE(4'b0000)
  ) lc40_16_29_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_67789),
    .in1(net_67790),
    .in2(net_67791_cascademuxed),
    .in3(net_67792),
    .lcout(net_63884),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_29_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_67835),
    .clk(net_67836),
    .in0(gnd),
    .in1(net_67802),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_63886),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011110000011100),
    .SEQ_MODE(4'b0000)
  ) lc40_16_29_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_67813),
    .in1(net_67814),
    .in2(net_67815_cascademuxed),
    .in3(net_67816),
    .lcout(net_63888),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_29_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_67825),
    .in1(gnd),
    .in2(net_67827_cascademuxed),
    .in3(gnd),
    .lcout(net_63890),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_16_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_64514),
    .clk(net_64515),
    .in0(gnd),
    .in1(net_64475),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_60528),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010100000110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_64480),
    .in1(net_64481),
    .in2(gnd),
    .in3(net_64483),
    .lcout(net_60529),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000110010),
    .SEQ_MODE(4'b0000)
  ) lc40_16_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_64486),
    .in1(gnd),
    .in2(net_64488_cascademuxed),
    .in3(gnd),
    .lcout(net_60530),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010100000001),
    .SEQ_MODE(4'b0000)
  ) lc40_16_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_64498),
    .in1(net_64499),
    .in2(net_64500_cascademuxed),
    .in3(net_64501),
    .lcout(net_60532),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_4_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_0 (
    .carryin(t450),
    .carryout(t452),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64838),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_1 (
    .carryin(t452),
    .carryout(net_64842),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_64845_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_2 (
    .carryin(net_64842),
    .carryout(net_64848),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64850),
    .in2(gnd),
    .in3(net_64852),
    .lcout(net_60934),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_3 (
    .carryin(net_64848),
    .carryout(net_64854),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64856),
    .in2(gnd),
    .in3(net_64858),
    .lcout(net_60935),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_4 (
    .carryin(net_64854),
    .carryout(net_64860),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64862),
    .in2(gnd),
    .in3(net_64864),
    .lcout(net_60936),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_5 (
    .carryin(net_64860),
    .carryout(net_64866),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64868),
    .in2(gnd),
    .in3(net_64870),
    .lcout(net_60937),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_6 (
    .carryin(net_64866),
    .carryout(net_64872),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64874),
    .in2(gnd),
    .in3(net_64876),
    .lcout(net_60938),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_5_7 (
    .carryin(net_64872),
    .carryout(net_64878),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_64880),
    .in2(gnd),
    .in3(net_64882),
    .lcout(net_60939),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_16_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_64962_cascademuxed),
    .in3(net_64963),
    .lcout(net_61055),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65341),
    .in1(net_65342),
    .in2(net_65343_cascademuxed),
    .in3(net_65344),
    .lcout(net_61426),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_9_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65375),
    .clk(net_65376),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_65350),
    .lcout(net_61427),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_16_9_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_65375),
    .clk(net_65376),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65355_cascademuxed),
    .in3(gnd),
    .lcout(net_61428),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65359),
    .in1(net_65360),
    .in2(net_65361_cascademuxed),
    .in3(net_65362),
    .lcout(net_61429),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_16_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_65367_cascademuxed),
    .in3(gnd),
    .lcout(net_61430),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_16_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_65371),
    .in1(net_65372),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_61431),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69576),
    .in0(net_69535),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65625),
    .ltout(),
    .sr(net_69577)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69698),
    .clk(net_69699),
    .in0(net_69670),
    .in1(net_69671),
    .in2(gnd),
    .in3(net_69673),
    .lcout(net_65750),
    .ltout(),
    .sr(net_69700)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000001000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69698),
    .clk(net_69699),
    .in0(gnd),
    .in1(net_69689),
    .in2(net_69690_cascademuxed),
    .in3(net_69691),
    .lcout(net_65753),
    .ltout(),
    .sr(net_69700)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69822),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69778),
    .lcout(net_65870),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69822),
    .in0(gnd),
    .in1(net_69788),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65872),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69822),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69796),
    .lcout(net_65873),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69822),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_69802),
    .lcout(net_65874),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110011111111),
    .SEQ_MODE(4'b0000)
  ) lc40_17_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_69805),
    .in1(net_69806),
    .in2(net_69807_cascademuxed),
    .in3(net_69808),
    .lcout(net_65875),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_69822),
    .in0(net_69817),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65877),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_69898),
    .in1(gnd),
    .in2(net_69900_cascademuxed),
    .in3(gnd),
    .lcout(net_65993),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100100011),
    .SEQ_MODE(4'b0000)
  ) lc40_17_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_69916),
    .in1(gnd),
    .in2(net_69918_cascademuxed),
    .in3(net_69919),
    .lcout(net_65996),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69944),
    .clk(net_69945),
    .in0(gnd),
    .in1(net_69923),
    .in2(net_69924_cascademuxed),
    .in3(net_69925),
    .lcout(net_65997),
    .ltout(),
    .sr(net_69946)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_16_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70068),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_70030),
    .lcout(net_66117),
    .ltout(),
    .sr(net_70069)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_17_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70065_cascademuxed),
    .in3(gnd),
    .lcout(net_66123),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70190),
    .clk(net_70191),
    .in0(gnd),
    .in1(net_70145),
    .in2(net_70146_cascademuxed),
    .in3(net_70147),
    .lcout(net_66239),
    .ltout(),
    .sr(net_70192)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_70150),
    .in1(net_70151),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_66240),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000010111000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70190),
    .clk(net_70191),
    .in0(net_70156),
    .in1(net_70157),
    .in2(net_70158_cascademuxed),
    .in3(gnd),
    .lcout(net_66241),
    .ltout(),
    .sr(net_70192)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001010100),
    .SEQ_MODE(4'b0000)
  ) lc40_17_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70175),
    .in2(net_70176_cascademuxed),
    .in3(gnd),
    .lcout(net_66244),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000110101),
    .SEQ_MODE(4'b0000)
  ) lc40_17_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_70186),
    .in1(net_70187),
    .in2(net_70188_cascademuxed),
    .in3(gnd),
    .lcout(net_66246),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70314),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70269_cascademuxed),
    .in3(gnd),
    .lcout(net_66362),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70314),
    .in0(gnd),
    .in1(net_70274),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_66363),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70314),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_70282),
    .lcout(net_66364),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70314),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_70288),
    .lcout(net_66365),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70314),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70293_cascademuxed),
    .in3(gnd),
    .lcout(net_66366),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70314),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70305_cascademuxed),
    .in3(gnd),
    .lcout(net_66368),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_70314),
    .in0(net_70309),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_66369),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_19_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70436),
    .clk(net_70437),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70398_cascademuxed),
    .in3(gnd),
    .lcout(net_66486),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101110111011),
    .SEQ_MODE(4'b0000)
  ) lc40_17_19_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_70414),
    .in1(net_70415),
    .in2(net_70416_cascademuxed),
    .in3(net_70417),
    .lcout(net_66489),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_19_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70436),
    .clk(net_70437),
    .in0(net_70420),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_66490),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101110111011),
    .SEQ_MODE(4'b0000)
  ) lc40_17_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_70426),
    .in1(net_70427),
    .in2(net_70428_cascademuxed),
    .in3(net_70429),
    .lcout(net_66491),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_70433),
    .in2(net_70434_cascademuxed),
    .in3(gnd),
    .lcout(net_66492),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_20_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70559),
    .clk(net_70560),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70515_cascademuxed),
    .in3(gnd),
    .lcout(net_66608),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111110110011),
    .SEQ_MODE(4'b0000)
  ) lc40_17_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_70519),
    .in1(net_70520),
    .in2(net_70521_cascademuxed),
    .in3(net_70522),
    .lcout(net_66609),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_20_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70559),
    .clk(net_70560),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_70528),
    .lcout(net_66610),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_20_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70559),
    .clk(net_70560),
    .in0(net_70543),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_66613),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_20_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_70549),
    .in1(net_70550),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_66614),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_21_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70682),
    .clk(net_70683),
    .in0(gnd),
    .in1(gnd),
    .in2(net_70668_cascademuxed),
    .in3(gnd),
    .lcout(net_66736),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_21_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_70682),
    .clk(net_70683),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_70675),
    .lcout(net_66737),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000011111111000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_29_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_71650),
    .in1(net_71651),
    .in2(net_71652_cascademuxed),
    .in3(net_71653),
    .lcout(net_67720),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000101000101010),
    .SEQ_MODE(4'b0000)
  ) lc40_17_29_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_71656),
    .in1(net_71657),
    .in2(net_71658_cascademuxed),
    .in3(net_71659),
    .lcout(net_67721),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010111101110),
    .SEQ_MODE(4'b0000)
  ) lc40_17_29_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_71662),
    .in1(net_71663),
    .in2(net_71664_cascademuxed),
    .in3(net_71665),
    .lcout(net_67722),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68714),
    .clk(net_68715),
    .in0(gnd),
    .in1(gnd),
    .in2(net_68670_cascademuxed),
    .in3(net_68671),
    .lcout(net_64763),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68714),
    .clk(net_68715),
    .in0(gnd),
    .in1(net_68675),
    .in2(gnd),
    .in3(net_68677),
    .lcout(net_64764),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68714),
    .clk(net_68715),
    .in0(net_68680),
    .in1(net_68681),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_64765),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68714),
    .clk(net_68715),
    .in0(gnd),
    .in1(net_68687),
    .in2(gnd),
    .in3(net_68689),
    .lcout(net_64766),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_68698),
    .in1(net_68699),
    .in2(gnd),
    .in3(net_68701),
    .lcout(net_64768),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68714),
    .clk(net_68715),
    .in0(gnd),
    .in1(net_68705),
    .in2(net_68706_cascademuxed),
    .in3(gnd),
    .lcout(net_64769),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68714),
    .clk(net_68715),
    .in0(gnd),
    .in1(net_68711),
    .in2(net_68712_cascademuxed),
    .in3(gnd),
    .lcout(net_64770),
    .ltout(),
    .sr(net_68716)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_17_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_68837),
    .clk(net_68838),
    .in0(gnd),
    .in1(net_68792),
    .in2(gnd),
    .in3(net_68794),
    .lcout(net_64886),
    .ltout(),
    .sr(net_68839)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b0000)
  ) lc40_17_6_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_68815),
    .in1(net_68816),
    .in2(net_68817_cascademuxed),
    .in3(gnd),
    .lcout(net_64890),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_17_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_68821),
    .in1(net_68822),
    .in2(net_68823_cascademuxed),
    .in3(net_68824),
    .lcout(net_64891),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_17_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_68833),
    .in1(net_68834),
    .in2(net_68835_cascademuxed),
    .in3(net_68836),
    .lcout(net_64893),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_17_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_69206),
    .clk(net_69207),
    .in0(net_69166),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_65256),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100010001),
    .SEQ_MODE(4'b0000)
  ) lc40_18_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_73132),
    .in1(net_73133),
    .in2(net_73134_cascademuxed),
    .in3(net_73135),
    .lcout(net_69212),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(net_73378),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69458),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(net_73396),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69461),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73407),
    .in0(net_73402),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69462),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(net_73484),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69578),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73492),
    .lcout(net_69579),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73497_cascademuxed),
    .in3(gnd),
    .lcout(net_69580),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000010101),
    .SEQ_MODE(4'b0000)
  ) lc40_18_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_73502),
    .in2(net_73503_cascademuxed),
    .in3(net_73504),
    .lcout(net_69581),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100110001),
    .SEQ_MODE(4'b0000)
  ) lc40_18_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_73507),
    .in1(gnd),
    .in2(net_73509_cascademuxed),
    .in3(net_73510),
    .lcout(net_69582),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(net_73514),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69583),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73522),
    .lcout(net_69584),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73530),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73527_cascademuxed),
    .in3(gnd),
    .lcout(net_69585),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011100100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_73652),
    .clk(net_73653),
    .in0(net_73606),
    .in1(net_73607),
    .in2(net_73608_cascademuxed),
    .in3(gnd),
    .lcout(net_69701),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000101000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_73652),
    .clk(net_73653),
    .in0(gnd),
    .in1(net_73613),
    .in2(net_73614_cascademuxed),
    .in3(net_73615),
    .lcout(net_69702),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000111),
    .SEQ_MODE(4'b0000)
  ) lc40_18_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_73618),
    .in1(net_73619),
    .in2(gnd),
    .in3(net_73621),
    .lcout(net_69703),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010100000011),
    .SEQ_MODE(4'b0000)
  ) lc40_18_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_73624),
    .in1(net_73625),
    .in2(gnd),
    .in3(net_73627),
    .lcout(net_69704),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_73652),
    .clk(net_73653),
    .in0(net_73630),
    .in1(gnd),
    .in2(net_73632_cascademuxed),
    .in3(net_73633),
    .lcout(net_69705),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000101000001100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_73652),
    .clk(net_73653),
    .in0(net_73636),
    .in1(net_73637),
    .in2(gnd),
    .in3(net_73639),
    .lcout(net_69706),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011000000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_73652),
    .clk(net_73653),
    .in0(net_73648),
    .in1(gnd),
    .in2(net_73650_cascademuxed),
    .in3(net_73651),
    .lcout(net_69708),
    .ltout(),
    .sr(net_73654)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73776),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73732),
    .lcout(net_69824),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73776),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73744),
    .lcout(net_69826),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73776),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73749_cascademuxed),
    .in3(gnd),
    .lcout(net_69827),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73776),
    .in0(net_73753),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69828),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73776),
    .in0(net_73759),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69829),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73776),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73767_cascademuxed),
    .in3(gnd),
    .lcout(net_69830),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73776),
    .in0(net_73771),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_69831),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_18_16_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_73899),
    .in0(gnd),
    .in1(net_73865),
    .in2(gnd),
    .in3(net_73867),
    .lcout(net_69949),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74022),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_73978),
    .lcout(net_70070),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74022),
    .in0(gnd),
    .in1(gnd),
    .in2(net_73983_cascademuxed),
    .in3(gnd),
    .lcout(net_70071),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74022),
    .in0(net_73987),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_70072),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74022),
    .in0(gnd),
    .in1(net_73994),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_70073),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74022),
    .in0(gnd),
    .in1(gnd),
    .in2(net_74001_cascademuxed),
    .in3(gnd),
    .lcout(net_70074),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010001100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_74005),
    .in1(net_74006),
    .in2(net_74007_cascademuxed),
    .in3(net_74008),
    .lcout(net_70075),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74022),
    .in0(gnd),
    .in1(gnd),
    .in2(net_74013_cascademuxed),
    .in3(gnd),
    .lcout(net_70076),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74022),
    .in0(gnd),
    .in1(net_74018),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_70077),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010101000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_74144),
    .clk(net_74145),
    .in0(gnd),
    .in1(net_74111),
    .in2(net_74112_cascademuxed),
    .in3(net_74113),
    .lcout(net_70195),
    .ltout(),
    .sr(net_74146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_74144),
    .clk(net_74145),
    .in0(net_74116),
    .in1(net_74117),
    .in2(gnd),
    .in3(net_74119),
    .lcout(net_70196),
    .ltout(),
    .sr(net_74146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100100011),
    .SEQ_MODE(4'b0000)
  ) lc40_18_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_74122),
    .in1(gnd),
    .in2(net_74124_cascademuxed),
    .in3(net_74125),
    .lcout(net_70197),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_74144),
    .clk(net_74145),
    .in0(net_74128),
    .in1(net_74129),
    .in2(gnd),
    .in3(net_74131),
    .lcout(net_70198),
    .ltout(),
    .sr(net_74146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110100001000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_74144),
    .clk(net_74145),
    .in0(net_74134),
    .in1(net_74135),
    .in2(gnd),
    .in3(net_74137),
    .lcout(net_70199),
    .ltout(),
    .sr(net_74146)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001100000101),
    .SEQ_MODE(4'b0000)
  ) lc40_18_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_74140),
    .in1(net_74141),
    .in2(gnd),
    .in3(net_74143),
    .lcout(net_70200),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_18_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_74267),
    .clk(net_74268),
    .in0(net_74263),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_70323),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_18_20_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_74391),
    .in0(gnd),
    .in1(net_74387),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_70446),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_18_5_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_72545),
    .clk(net_72546),
    .in0(gnd),
    .in1(net_72530),
    .in2(gnd),
    .in3(net_72532),
    .lcout(net_68599),
    .ltout(),
    .sr(net_72547)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_18_5_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_72541),
    .in1(gnd),
    .in2(gnd),
    .in3(net_72544),
    .lcout(net_68601),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_72622),
    .in1(gnd),
    .in2(net_72624_cascademuxed),
    .in3(net_72625),
    .lcout(net_68717),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_6_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_72628),
    .in1(net_72629),
    .in2(net_72630_cascademuxed),
    .in3(net_72631),
    .lcout(net_68718),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_18_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72635),
    .in2(gnd),
    .in3(net_72637),
    .lcout(net_68719),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001010101010101),
    .SEQ_MODE(4'b0000)
  ) lc40_18_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_72652),
    .in1(net_72653),
    .in2(net_72654_cascademuxed),
    .in3(net_72655),
    .lcout(net_68722),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_18_6_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_72659),
    .in2(net_72660_cascademuxed),
    .in3(net_72661),
    .lcout(net_68723),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_18_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_72668),
    .clk(net_72669),
    .in0(net_72664),
    .in1(gnd),
    .in2(net_72666_cascademuxed),
    .in3(gnd),
    .lcout(net_68724),
    .ltout(),
    .sr(net_72670)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100110011001100),
    .SEQ_MODE(4'b0000)
  ) lc40_1_30_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_11052),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_20_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_80146),
    .in2(net_80147_cascademuxed),
    .in3(net_80148),
    .lcout(net_76651),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_20_10_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80163),
    .in1(net_80164),
    .in2(net_80165_cascademuxed),
    .in3(net_80166),
    .lcout(net_76654),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100111111001010),
    .SEQ_MODE(4'b0000)
  ) lc40_20_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80175),
    .in1(net_80176),
    .in2(net_80177_cascademuxed),
    .in3(net_80178),
    .lcout(net_76656),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80191),
    .clk(net_80192),
    .in0(net_80187),
    .in1(gnd),
    .in2(net_80189_cascademuxed),
    .in3(gnd),
    .lcout(net_76658),
    .ltout(),
    .sr(net_80193)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80315),
    .in0(gnd),
    .in1(gnd),
    .in2(net_80300_cascademuxed),
    .in3(gnd),
    .lcout(net_76758),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000101010001),
    .SEQ_MODE(4'b0000)
  ) lc40_20_12_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_80392),
    .in2(net_80393_cascademuxed),
    .in3(net_80394),
    .lcout(net_76855),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110100001000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80437),
    .clk(net_80438),
    .in0(net_80397),
    .in1(net_80398),
    .in2(gnd),
    .in3(net_80400),
    .lcout(net_76856),
    .ltout(),
    .sr(net_80439)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000101000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80437),
    .clk(net_80438),
    .in0(gnd),
    .in1(net_80404),
    .in2(net_80405_cascademuxed),
    .in3(net_80406),
    .lcout(net_76857),
    .ltout(),
    .sr(net_80439)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110100001000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80437),
    .clk(net_80438),
    .in0(net_80409),
    .in1(net_80410),
    .in2(gnd),
    .in3(net_80412),
    .lcout(net_76858),
    .ltout(),
    .sr(net_80439)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000010011),
    .SEQ_MODE(4'b0000)
  ) lc40_20_12_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80415),
    .in1(gnd),
    .in2(net_80417_cascademuxed),
    .in3(net_80418),
    .lcout(net_76859),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80437),
    .clk(net_80438),
    .in0(net_80421),
    .in1(net_80422),
    .in2(gnd),
    .in3(net_80424),
    .lcout(net_76860),
    .ltout(),
    .sr(net_80439)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000101000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_12_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80437),
    .clk(net_80438),
    .in0(gnd),
    .in1(net_80428),
    .in2(net_80429_cascademuxed),
    .in3(net_80430),
    .lcout(net_76861),
    .ltout(),
    .sr(net_80439)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001100010001),
    .SEQ_MODE(4'b0000)
  ) lc40_20_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80433),
    .in1(gnd),
    .in2(net_80435_cascademuxed),
    .in3(net_80436),
    .lcout(net_76862),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100001011),
    .SEQ_MODE(4'b0000)
  ) lc40_20_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80514),
    .in1(net_80515),
    .in2(net_80516_cascademuxed),
    .in3(net_80517),
    .lcout(net_76957),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80560),
    .clk(net_80561),
    .in0(gnd),
    .in1(net_80521),
    .in2(net_80522_cascademuxed),
    .in3(net_80523),
    .lcout(net_76958),
    .ltout(),
    .sr(net_80562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011000100100000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80560),
    .clk(net_80561),
    .in0(net_80526),
    .in1(gnd),
    .in2(net_80528_cascademuxed),
    .in3(net_80529),
    .lcout(net_76959),
    .ltout(),
    .sr(net_80562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80560),
    .clk(net_80561),
    .in0(net_80532),
    .in1(net_80533),
    .in2(gnd),
    .in3(net_80535),
    .lcout(net_76960),
    .ltout(),
    .sr(net_80562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011001010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80560),
    .clk(net_80561),
    .in0(net_80538),
    .in1(net_80539),
    .in2(net_80540_cascademuxed),
    .in3(gnd),
    .lcout(net_76961),
    .ltout(),
    .sr(net_80562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80560),
    .clk(net_80561),
    .in0(net_80544),
    .in1(net_80545),
    .in2(gnd),
    .in3(net_80547),
    .lcout(net_76962),
    .ltout(),
    .sr(net_80562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011100100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80560),
    .clk(net_80561),
    .in0(net_80550),
    .in1(net_80551),
    .in2(net_80552_cascademuxed),
    .in3(gnd),
    .lcout(net_76963),
    .ltout(),
    .sr(net_80562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011100010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80560),
    .clk(net_80561),
    .in0(net_80556),
    .in1(net_80557),
    .in2(net_80558_cascademuxed),
    .in3(gnd),
    .lcout(net_76964),
    .ltout(),
    .sr(net_80562)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000111),
    .SEQ_MODE(4'b0000)
  ) lc40_20_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80637),
    .in1(net_80638),
    .in2(net_80639_cascademuxed),
    .in3(gnd),
    .lcout(net_77059),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80684),
    .in0(gnd),
    .in1(net_80644),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_77060),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80684),
    .in0(net_80649),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_77061),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000101000101),
    .SEQ_MODE(4'b0000)
  ) lc40_20_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80655),
    .in1(net_80656),
    .in2(net_80657_cascademuxed),
    .in3(net_80658),
    .lcout(net_77062),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80684),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_80664),
    .lcout(net_77063),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000010011),
    .SEQ_MODE(4'b0000)
  ) lc40_20_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80667),
    .in1(gnd),
    .in2(net_80669_cascademuxed),
    .in3(net_80670),
    .lcout(net_77064),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000111),
    .SEQ_MODE(4'b0000)
  ) lc40_20_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80673),
    .in1(net_80674),
    .in2(gnd),
    .in3(net_80676),
    .lcout(net_77065),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000101000101),
    .SEQ_MODE(4'b0000)
  ) lc40_20_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80679),
    .in1(net_80680),
    .in2(net_80681_cascademuxed),
    .in3(net_80682),
    .lcout(net_77066),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000110101),
    .SEQ_MODE(4'b0000)
  ) lc40_20_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80760),
    .in1(net_80761),
    .in2(net_80762_cascademuxed),
    .in3(gnd),
    .lcout(net_77161),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80806),
    .clk(net_80807),
    .in0(gnd),
    .in1(net_80767),
    .in2(net_80768_cascademuxed),
    .in3(net_80769),
    .lcout(net_77162),
    .ltout(),
    .sr(net_80808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011000000100010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80806),
    .clk(net_80807),
    .in0(net_80772),
    .in1(gnd),
    .in2(net_80774_cascademuxed),
    .in3(net_80775),
    .lcout(net_77163),
    .ltout(),
    .sr(net_80808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80806),
    .clk(net_80807),
    .in0(net_80778),
    .in1(net_80779),
    .in2(net_80780_cascademuxed),
    .in3(gnd),
    .lcout(net_77164),
    .ltout(),
    .sr(net_80808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000101000001100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80806),
    .clk(net_80807),
    .in0(net_80784),
    .in1(net_80785),
    .in2(gnd),
    .in3(net_80787),
    .lcout(net_77165),
    .ltout(),
    .sr(net_80808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80806),
    .clk(net_80807),
    .in0(net_80790),
    .in1(net_80791),
    .in2(gnd),
    .in3(net_80793),
    .lcout(net_77166),
    .ltout(),
    .sr(net_80808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80806),
    .clk(net_80807),
    .in0(gnd),
    .in1(net_80797),
    .in2(net_80798_cascademuxed),
    .in3(net_80799),
    .lcout(net_77167),
    .ltout(),
    .sr(net_80808)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011000100100000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80806),
    .clk(net_80807),
    .in0(net_80802),
    .in1(gnd),
    .in2(net_80804_cascademuxed),
    .in3(net_80805),
    .lcout(net_77168),
    .ltout(),
    .sr(net_80808)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_20_16_0 (
    .carryin(t630),
    .carryout(net_80882),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_80884),
    .in2(net_80885_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_20_16_1 (
    .carryin(net_80882),
    .carryout(net_80888),
    .ce(),
    .clk(net_80930),
    .in0(gnd),
    .in1(net_80890),
    .in2(gnd),
    .in3(net_80892),
    .lcout(net_77264),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_20_16_2 (
    .carryin(net_80888),
    .carryout(net_80894),
    .ce(),
    .clk(net_80930),
    .in0(gnd),
    .in1(gnd),
    .in2(net_80897_cascademuxed),
    .in3(net_80898),
    .lcout(net_77265),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_20_16_3 (
    .carryin(net_80894),
    .carryout(net_80900),
    .ce(),
    .clk(net_80930),
    .in0(gnd),
    .in1(net_80902),
    .in2(gnd),
    .in3(net_80904),
    .lcout(net_77266),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_20_16_4 (
    .carryin(net_80900),
    .carryout(net_80906),
    .ce(),
    .clk(net_80930),
    .in0(gnd),
    .in1(net_80908),
    .in2(gnd),
    .in3(net_80910),
    .lcout(net_77267),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_20_16_5 (
    .carryin(net_80906),
    .carryout(net_80912),
    .ce(),
    .clk(net_80930),
    .in0(gnd),
    .in1(gnd),
    .in2(net_80915_cascademuxed),
    .in3(net_80916),
    .lcout(net_77268),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_20_16_6 (
    .carryin(net_80912),
    .carryout(net_80918),
    .ce(),
    .clk(net_80930),
    .in0(gnd),
    .in1(net_80920),
    .in2(gnd),
    .in3(net_80922),
    .lcout(net_77269),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_20_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_80930),
    .in0(gnd),
    .in1(net_80926),
    .in2(gnd),
    .in3(net_80928),
    .lcout(net_77270),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000110000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_20_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_81006),
    .in1(net_81007),
    .in2(net_81008_cascademuxed),
    .in3(net_81009),
    .lcout(net_77365),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010001100100000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_81052),
    .clk(net_81053),
    .in0(net_81012),
    .in1(gnd),
    .in2(net_81014_cascademuxed),
    .in3(net_81015),
    .lcout(net_77366),
    .ltout(),
    .sr(net_81054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000010000100001),
    .SEQ_MODE(4'b0000)
  ) lc40_20_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_81018),
    .in1(net_81019),
    .in2(net_81020_cascademuxed),
    .in3(net_81021),
    .lcout(net_77367),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110100001000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_81052),
    .clk(net_81053),
    .in0(net_81024),
    .in1(net_81025),
    .in2(gnd),
    .in3(net_81027),
    .lcout(net_77368),
    .ltout(),
    .sr(net_81054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100010000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_20_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_81030),
    .in1(net_81031),
    .in2(net_81032_cascademuxed),
    .in3(net_81033),
    .lcout(net_77369),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010001100100000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_81052),
    .clk(net_81053),
    .in0(net_81036),
    .in1(gnd),
    .in2(net_81038_cascademuxed),
    .in3(net_81039),
    .lcout(net_77370),
    .ltout(),
    .sr(net_81054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000101000101),
    .SEQ_MODE(4'b0000)
  ) lc40_20_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_81043),
    .in2(net_81044_cascademuxed),
    .in3(net_81045),
    .lcout(net_77371),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_81052),
    .clk(net_81053),
    .in0(net_81048),
    .in1(gnd),
    .in2(net_81050_cascademuxed),
    .in3(net_81051),
    .lcout(net_77372),
    .ltout(),
    .sr(net_81054)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_81175),
    .clk(net_81176),
    .in0(net_81135),
    .in1(net_81136),
    .in2(gnd),
    .in3(net_81138),
    .lcout(net_77468),
    .ltout(),
    .sr(net_81177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_81175),
    .clk(net_81176),
    .in0(gnd),
    .in1(net_81148),
    .in2(net_81149_cascademuxed),
    .in3(net_81150),
    .lcout(net_77470),
    .ltout(),
    .sr(net_81177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011100100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_81175),
    .clk(net_81176),
    .in0(net_81153),
    .in1(net_81154),
    .in2(net_81155_cascademuxed),
    .in3(gnd),
    .lcout(net_77471),
    .ltout(),
    .sr(net_81177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000010100010),
    .SEQ_MODE(4'b0000)
  ) lc40_20_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_81159),
    .in1(net_81160),
    .in2(net_81161_cascademuxed),
    .in3(net_81162),
    .lcout(net_77472),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000001000100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_81175),
    .clk(net_81176),
    .in0(gnd),
    .in1(net_81172),
    .in2(net_81173_cascademuxed),
    .in3(net_81174),
    .lcout(net_77474),
    .ltout(),
    .sr(net_81177)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_20_19_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_81299),
    .in0(gnd),
    .in1(net_81289),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_77575),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_20_19_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_81299),
    .in0(net_81294),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_77576),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_20_6_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_79653),
    .in1(net_79654),
    .in2(net_79655_cascademuxed),
    .in3(net_79656),
    .lcout(net_76243),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_20_6_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_79667_cascademuxed),
    .in3(net_79668),
    .lcout(net_76245),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79699),
    .clk(net_79700),
    .in0(gnd),
    .in1(gnd),
    .in2(net_79685_cascademuxed),
    .in3(net_79686),
    .lcout(net_76248),
    .ltout(),
    .sr(net_79701)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_20_6_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_79699),
    .clk(net_79700),
    .in0(gnd),
    .in1(gnd),
    .in2(net_79697_cascademuxed),
    .in3(gnd),
    .lcout(net_76250),
    .ltout(),
    .sr(net_79701)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100011),
    .SEQ_MODE(4'b0000)
  ) lc40_20_7_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_79776),
    .in1(gnd),
    .in2(net_79778_cascademuxed),
    .in3(gnd),
    .lcout(net_76345),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001100000010),
    .SEQ_MODE(4'b0000)
  ) lc40_20_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_80022),
    .in1(gnd),
    .in2(gnd),
    .in3(net_80025),
    .lcout(net_76549),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_20_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_80068),
    .clk(net_80069),
    .in0(net_80028),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_76550),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_20_9_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_80053),
    .in2(gnd),
    .in3(net_80055),
    .lcout(net_76554),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_21_10_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_83976),
    .in1(gnd),
    .in2(net_83978_cascademuxed),
    .in3(gnd),
    .lcout(net_80071),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84022),
    .clk(net_84023),
    .in0(net_83982),
    .in1(gnd),
    .in2(gnd),
    .in3(net_83985),
    .lcout(net_80072),
    .ltout(),
    .sr(net_84024)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84022),
    .clk(net_84023),
    .in0(gnd),
    .in1(net_84001),
    .in2(net_84002_cascademuxed),
    .in3(gnd),
    .lcout(net_80075),
    .ltout(),
    .sr(net_84024)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111100001110),
    .SEQ_MODE(4'b0000)
  ) lc40_21_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84006),
    .in1(net_84007),
    .in2(gnd),
    .in3(net_84009),
    .lcout(net_80076),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84269),
    .in0(gnd),
    .in1(net_84235),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_80319),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000110101),
    .SEQ_MODE(4'b0000)
  ) lc40_21_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84252),
    .in1(net_84253),
    .in2(net_84254_cascademuxed),
    .in3(net_84255),
    .lcout(net_80322),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84269),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_84267),
    .lcout(net_80324),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000011001010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_13_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84391),
    .clk(net_84392),
    .in0(net_84345),
    .in1(net_84346),
    .in2(net_84347_cascademuxed),
    .in3(gnd),
    .lcout(net_80440),
    .ltout(),
    .sr(net_84393)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001010011),
    .SEQ_MODE(4'b0000)
  ) lc40_21_13_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84351),
    .in1(net_84352),
    .in2(net_84353_cascademuxed),
    .in3(gnd),
    .lcout(net_80441),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100100011),
    .SEQ_MODE(4'b0000)
  ) lc40_21_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84357),
    .in1(net_84358),
    .in2(net_84359_cascademuxed),
    .in3(net_84360),
    .lcout(net_80442),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_13_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84391),
    .clk(net_84392),
    .in0(net_84363),
    .in1(net_84364),
    .in2(gnd),
    .in3(net_84366),
    .lcout(net_80443),
    .ltout(),
    .sr(net_84393)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_13_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84391),
    .clk(net_84392),
    .in0(net_84369),
    .in1(net_84370),
    .in2(net_84371_cascademuxed),
    .in3(gnd),
    .lcout(net_80444),
    .ltout(),
    .sr(net_84393)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84391),
    .clk(net_84392),
    .in0(net_84381),
    .in1(net_84382),
    .in2(net_84383_cascademuxed),
    .in3(gnd),
    .lcout(net_80446),
    .ltout(),
    .sr(net_84393)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000110000001010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84391),
    .clk(net_84392),
    .in0(net_84387),
    .in1(net_84388),
    .in2(gnd),
    .in3(net_84390),
    .lcout(net_80447),
    .ltout(),
    .sr(net_84393)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_21_14_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84468),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_80563),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110111011110000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_14_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84514),
    .clk(net_84515),
    .in0(net_84474),
    .in1(net_84475),
    .in2(net_84476_cascademuxed),
    .in3(net_84477),
    .lcout(net_80564),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101111001000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84514),
    .clk(net_84515),
    .in0(net_84480),
    .in1(net_84481),
    .in2(net_84482_cascademuxed),
    .in3(net_84483),
    .lcout(net_80565),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101011001010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84514),
    .clk(net_84515),
    .in0(net_84486),
    .in1(net_84487),
    .in2(net_84488_cascademuxed),
    .in3(net_84489),
    .lcout(net_80566),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110010101100),
    .SEQ_MODE(4'b1000)
  ) lc40_21_14_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84514),
    .clk(net_84515),
    .in0(net_84492),
    .in1(net_84493),
    .in2(net_84494_cascademuxed),
    .in3(net_84495),
    .lcout(net_80567),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111101111001000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_14_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84514),
    .clk(net_84515),
    .in0(net_84498),
    .in1(net_84499),
    .in2(net_84500_cascademuxed),
    .in3(net_84501),
    .lcout(net_80568),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110110101000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_14_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84514),
    .clk(net_84515),
    .in0(net_84504),
    .in1(net_84505),
    .in2(net_84506_cascademuxed),
    .in3(net_84507),
    .lcout(net_80569),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111110010101010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_14_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84514),
    .clk(net_84515),
    .in0(net_84510),
    .in1(net_84511),
    .in2(net_84512_cascademuxed),
    .in3(net_84513),
    .lcout(net_80570),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011001011111110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_15_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84637),
    .clk(net_84638),
    .in0(net_84591),
    .in1(net_84592),
    .in2(net_84593_cascademuxed),
    .in3(net_84594),
    .lcout(net_80686),
    .ltout(),
    .sr(net_84639)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100110001),
    .SEQ_MODE(4'b0000)
  ) lc40_21_15_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84597),
    .in1(net_84598),
    .in2(net_84599_cascademuxed),
    .in3(net_84600),
    .lcout(net_80687),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001110010),
    .SEQ_MODE(4'b0000)
  ) lc40_21_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84603),
    .in1(net_84604),
    .in2(net_84605_cascademuxed),
    .in3(gnd),
    .lcout(net_80688),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001100000101),
    .SEQ_MODE(4'b0000)
  ) lc40_21_15_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84609),
    .in1(net_84610),
    .in2(gnd),
    .in3(net_84612),
    .lcout(net_80689),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000010011),
    .SEQ_MODE(4'b0000)
  ) lc40_21_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84615),
    .in1(gnd),
    .in2(net_84617_cascademuxed),
    .in3(net_84618),
    .lcout(net_80690),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001100010001),
    .SEQ_MODE(4'b0000)
  ) lc40_21_15_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84621),
    .in1(net_84622),
    .in2(net_84623_cascademuxed),
    .in3(net_84624),
    .lcout(net_80691),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010101000000),
    .SEQ_MODE(4'b0000)
  ) lc40_21_15_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84627),
    .in1(net_84628),
    .in2(net_84629_cascademuxed),
    .in3(net_84630),
    .lcout(net_80692),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000110100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_21_15_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84633),
    .in1(net_84634),
    .in2(net_84635_cascademuxed),
    .in3(net_84636),
    .lcout(net_80693),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_21_16_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84732),
    .in1(net_84733),
    .in2(net_84734_cascademuxed),
    .in3(net_84735),
    .lcout(net_80812),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_21_16_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_84739),
    .in2(gnd),
    .in3(net_84741),
    .lcout(net_80813),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_16_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_84760),
    .clk(net_84761),
    .in0(net_84750),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_80815),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000001001000001),
    .SEQ_MODE(4'b0000)
  ) lc40_21_17_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84837),
    .in1(net_84838),
    .in2(net_84839_cascademuxed),
    .in3(net_84840),
    .lcout(net_80932),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000001001000001),
    .SEQ_MODE(4'b0000)
  ) lc40_21_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84843),
    .in1(net_84844),
    .in2(net_84845_cascademuxed),
    .in3(net_84846),
    .lcout(net_80933),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000001001000001),
    .SEQ_MODE(4'b0000)
  ) lc40_21_17_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84849),
    .in1(net_84850),
    .in2(net_84851_cascademuxed),
    .in3(net_84852),
    .lcout(net_80934),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_17_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84884),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_84858),
    .lcout(net_80935),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_17_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84884),
    .in0(gnd),
    .in1(gnd),
    .in2(net_84863_cascademuxed),
    .in3(gnd),
    .lcout(net_80936),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84884),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_84870),
    .lcout(net_80937),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_17_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84884),
    .in0(net_84873),
    .in1(net_84874),
    .in2(net_84875_cascademuxed),
    .in3(net_84876),
    .lcout(net_80938),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_84884),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_84882),
    .lcout(net_80939),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_85006),
    .clk(net_85007),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_84963),
    .lcout(net_81055),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_21_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_85006),
    .clk(net_85007),
    .in0(net_84966),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_81056),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100001101),
    .SEQ_MODE(4'b0000)
  ) lc40_21_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84972),
    .in1(net_84973),
    .in2(gnd),
    .in3(net_84975),
    .lcout(net_81057),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_18_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_85006),
    .clk(net_85007),
    .in0(gnd),
    .in1(gnd),
    .in2(net_84980_cascademuxed),
    .in3(gnd),
    .lcout(net_81058),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010100000011),
    .SEQ_MODE(4'b0000)
  ) lc40_21_18_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84984),
    .in1(net_84985),
    .in2(gnd),
    .in3(net_84987),
    .lcout(net_81059),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100010000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_21_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84990),
    .in1(net_84991),
    .in2(net_84992_cascademuxed),
    .in3(net_84993),
    .lcout(net_81060),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010100000011),
    .SEQ_MODE(4'b0000)
  ) lc40_21_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_84996),
    .in1(net_84997),
    .in2(gnd),
    .in3(net_84999),
    .lcout(net_81061),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000110100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_21_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_85002),
    .in1(net_85003),
    .in2(net_85004_cascademuxed),
    .in3(net_85005),
    .lcout(net_81062),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_19_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_85129),
    .clk(net_85130),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_85098),
    .lcout(net_81180),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_21_19_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_85129),
    .clk(net_85130),
    .in0(gnd),
    .in1(gnd),
    .in2(net_85103_cascademuxed),
    .in3(gnd),
    .lcout(net_81181),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000001000101),
    .SEQ_MODE(4'b0000)
  ) lc40_21_6_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_83503),
    .in2(net_83504_cascademuxed),
    .in3(net_83505),
    .lcout(net_79582),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_21_6_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_83514),
    .in1(net_83515),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_79584),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_21_9_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_83899),
    .clk(net_83900),
    .in0(gnd),
    .in1(net_83854),
    .in2(net_83855_cascademuxed),
    .in3(gnd),
    .lcout(net_79948),
    .ltout(),
    .sr(net_83901)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001010100),
    .SEQ_MODE(4'b0000)
  ) lc40_21_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_83866),
    .in2(net_83867_cascademuxed),
    .in3(gnd),
    .lcout(net_79950),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111000000010),
    .SEQ_MODE(4'b0000)
  ) lc40_21_9_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_83889),
    .in1(net_83890),
    .in2(gnd),
    .in3(net_83892),
    .lcout(net_79954),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_13_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_88223),
    .in0(gnd),
    .in1(gnd),
    .in2(net_88190_cascademuxed),
    .in3(gnd),
    .lcout(net_84273),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_88223),
    .in0(gnd),
    .in1(gnd),
    .in2(net_88208_cascademuxed),
    .in3(gnd),
    .lcout(net_84276),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100010001010000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_14_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_88345),
    .clk(net_88346),
    .in0(gnd),
    .in1(net_88318),
    .in2(net_88319_cascademuxed),
    .in3(net_88320),
    .lcout(net_84397),
    .ltout(),
    .sr(net_88347)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_15_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_88469),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_88437),
    .lcout(net_84519),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_15_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_88469),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_88449),
    .lcout(net_84521),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_22_16_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_88591),
    .clk(net_88592),
    .in0(gnd),
    .in1(net_88588),
    .in2(gnd),
    .in3(net_88590),
    .lcout(net_84647),
    .ltout(),
    .sr(net_88593)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_22_17_0 (
    .carryin(t735),
    .carryout(net_88667),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_88669),
    .in2(net_88670_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_22_17_1 (
    .carryin(net_88667),
    .carryout(net_88673),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_88676_cascademuxed),
    .in3(net_88677),
    .lcout(net_84764),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_22_17_2 (
    .carryin(net_88673),
    .carryout(net_88679),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_88681),
    .in2(gnd),
    .in3(net_88683),
    .lcout(net_84765),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_22_17_3 (
    .carryin(net_88679),
    .carryout(net_88685),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_88687),
    .in2(gnd),
    .in3(net_88689),
    .lcout(net_84766),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_22_17_4 (
    .carryin(net_88685),
    .carryout(net_88691),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_88693),
    .in2(gnd),
    .in3(net_88695),
    .lcout(net_84767),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_22_17_5 (
    .carryin(net_88691),
    .carryout(net_88697),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_88699),
    .in2(gnd),
    .in3(net_88701),
    .lcout(net_84768),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_22_17_6 (
    .carryin(net_88697),
    .carryout(net_88703),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_88705),
    .in2(gnd),
    .in3(net_88707),
    .lcout(net_84769),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_22_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_88712_cascademuxed),
    .in3(net_88713),
    .lcout(net_84770),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_22_9_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_87730),
    .clk(net_87731),
    .in0(gnd),
    .in1(gnd),
    .in2(net_87692_cascademuxed),
    .in3(gnd),
    .lcout(net_83780),
    .ltout(),
    .sr(net_87732)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_23_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_23_9_0 (
    .carryin(t753),
    .carryout(t755),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_91516),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_23_9_1 (
    .carryin(t755),
    .carryout(net_91520),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_91522),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_23_9_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_91561),
    .clk(net_91562),
    .in0(gnd),
    .in1(gnd),
    .in2(net_91529_cascademuxed),
    .in3(net_91530),
    .lcout(net_87612),
    .ltout(),
    .sr(net_91563)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_23_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_91557),
    .in1(net_91558),
    .in2(gnd),
    .in3(net_91560),
    .lcout(net_87617),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_2_19_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_13558),
    .in1(net_13559),
    .in2(net_13560_cascademuxed),
    .in3(net_13561),
    .lcout(net_9360),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_8_0 (
    .carryin(t0),
    .carryout(t2),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_12206),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_8_1 (
    .carryin(t2),
    .carryout(net_12210),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12213_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_8_2 (
    .carryin(net_12210),
    .carryout(net_12216),
    .ce(),
    .clk(net_12252),
    .in0(gnd),
    .in1(net_12218),
    .in2(gnd),
    .in3(net_12220),
    .lcout(net_7745),
    .ltout(),
    .sr(net_12253)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_8_3 (
    .carryin(net_12216),
    .carryout(net_12222),
    .ce(),
    .clk(net_12252),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12225_cascademuxed),
    .in3(net_12226),
    .lcout(net_7746),
    .ltout(),
    .sr(net_12253)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_8_4 (
    .carryin(net_12222),
    .carryout(net_12228),
    .ce(),
    .clk(net_12252),
    .in0(gnd),
    .in1(gnd),
    .in2(net_12231_cascademuxed),
    .in3(net_12232),
    .lcout(net_7747),
    .ltout(),
    .sr(net_12253)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_2_8_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_12252),
    .in0(gnd),
    .in1(net_12236),
    .in2(gnd),
    .in3(net_12238),
    .lcout(net_7748),
    .ltout(),
    .sr(net_12253)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000100000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_8_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12241),
    .in1(net_12242),
    .in2(net_12243_cascademuxed),
    .in3(net_12244),
    .lcout(net_7749),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_2_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_12247),
    .in1(net_12248),
    .in2(net_12249_cascademuxed),
    .in3(gnd),
    .lcout(net_7750),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_12_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_13_0 (
    .carryin(t8),
    .carryout(t10),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_16652),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_13_1 (
    .carryin(t10),
    .carryout(net_16656),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16659_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_2 (
    .carryin(net_16656),
    .carryout(net_16662),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(gnd),
    .in2(net_16665_cascademuxed),
    .in3(net_16666),
    .lcout(net_12748),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_3 (
    .carryin(net_16662),
    .carryout(net_16668),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16670),
    .in2(gnd),
    .in3(net_16672),
    .lcout(net_12749),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_4 (
    .carryin(net_16668),
    .carryout(net_16674),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16676),
    .in2(gnd),
    .in3(net_16678),
    .lcout(net_12750),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_16698),
    .in0(gnd),
    .in1(net_16682),
    .in2(gnd),
    .in3(net_16684),
    .lcout(net_12751),
    .ltout(),
    .sr(net_16699)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0100000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_13_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_16687),
    .in1(net_16688),
    .in2(net_16689_cascademuxed),
    .in3(net_16690),
    .lcout(net_12752),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_13_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_16693),
    .in1(net_16694),
    .in2(net_16695_cascademuxed),
    .in3(gnd),
    .lcout(net_12753),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_3_14_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_16820),
    .clk(net_16821),
    .in0(net_16786),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12871),
    .ltout(),
    .sr(net_16822)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_17_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_18_0 (
    .carryin(t11),
    .carryout(t13),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_17267),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_3_18_1 (
    .carryin(t13),
    .carryout(net_17271),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_17273),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_2 (
    .carryin(net_17271),
    .carryout(net_17277),
    .ce(),
    .clk(net_17313),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17280_cascademuxed),
    .in3(net_17281),
    .lcout(net_13363),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_3 (
    .carryin(net_17277),
    .carryout(net_17283),
    .ce(),
    .clk(net_17313),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17286_cascademuxed),
    .in3(net_17287),
    .lcout(net_13364),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_4 (
    .carryin(net_17283),
    .carryout(net_17289),
    .ce(),
    .clk(net_17313),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17292_cascademuxed),
    .in3(net_17293),
    .lcout(net_13365),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_5 (
    .carryin(net_17289),
    .carryout(net_17295),
    .ce(),
    .clk(net_17313),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17298_cascademuxed),
    .in3(net_17299),
    .lcout(net_13366),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_6 (
    .carryin(net_17295),
    .carryout(net_17301),
    .ce(),
    .clk(net_17313),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17304_cascademuxed),
    .in3(net_17305),
    .lcout(net_13367),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_18_7 (
    .carryin(net_17301),
    .carryout(net_17307),
    .ce(),
    .clk(net_17313),
    .in0(gnd),
    .in1(net_17309),
    .in2(gnd),
    .in3(net_17311),
    .lcout(net_13368),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_0 (
    .carryin(net_17351),
    .carryout(net_17388),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(net_17390),
    .in2(gnd),
    .in3(net_17392),
    .lcout(net_13484),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_1 (
    .carryin(net_17388),
    .carryout(net_17394),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17397_cascademuxed),
    .in3(net_17398),
    .lcout(net_13485),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_2 (
    .carryin(net_17394),
    .carryout(net_17400),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(net_17402),
    .in2(gnd),
    .in3(net_17404),
    .lcout(net_13486),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_3 (
    .carryin(net_17400),
    .carryout(net_17406),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(net_17408),
    .in2(gnd),
    .in3(net_17410),
    .lcout(net_13487),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_4 (
    .carryin(net_17406),
    .carryout(net_17412),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17415_cascademuxed),
    .in3(net_17416),
    .lcout(net_13488),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_5 (
    .carryin(net_17412),
    .carryout(net_17418),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17421_cascademuxed),
    .in3(net_17422),
    .lcout(net_13489),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_6 (
    .carryin(net_17418),
    .carryout(net_17424),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17427_cascademuxed),
    .in3(net_17428),
    .lcout(net_13490),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_19_7 (
    .carryin(net_17424),
    .carryout(net_17430),
    .ce(),
    .clk(net_17436),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17433_cascademuxed),
    .in3(net_17434),
    .lcout(net_13491),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_0 (
    .carryin(net_17474),
    .carryout(net_17511),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17514_cascademuxed),
    .in3(net_17515),
    .lcout(net_13607),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_1 (
    .carryin(net_17511),
    .carryout(net_17517),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(net_17519),
    .in2(gnd),
    .in3(net_17521),
    .lcout(net_13608),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_2 (
    .carryin(net_17517),
    .carryout(net_17523),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17526_cascademuxed),
    .in3(net_17527),
    .lcout(net_13609),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_3 (
    .carryin(net_17523),
    .carryout(net_17529),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(net_17531),
    .in2(gnd),
    .in3(net_17533),
    .lcout(net_13610),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_4 (
    .carryin(net_17529),
    .carryout(net_17535),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(net_17537),
    .in2(gnd),
    .in3(net_17539),
    .lcout(net_13611),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_5 (
    .carryin(net_17535),
    .carryout(net_17541),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(gnd),
    .in2(net_17544_cascademuxed),
    .in3(net_17545),
    .lcout(net_13612),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_6 (
    .carryin(net_17541),
    .carryout(net_17547),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(net_17549),
    .in2(gnd),
    .in3(net_17551),
    .lcout(net_13613),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_20_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_17559),
    .in0(gnd),
    .in1(net_17555),
    .in2(gnd),
    .in3(net_17557),
    .lcout(net_13614),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_3_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_15960),
    .in0(net_15955),
    .in1(gnd),
    .in2(gnd),
    .in3(net_15958),
    .lcout(net_12015),
    .ltout(),
    .sr(net_15961)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_3_8_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_16082),
    .clk(net_16083),
    .in0(gnd),
    .in1(net_16061),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_12135),
    .ltout(),
    .sr(net_16084)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20406),
    .in0(net_20371),
    .in1(gnd),
    .in2(gnd),
    .in3(net_20374),
    .lcout(net_16456),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_13_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_20529),
    .in0(gnd),
    .in1(net_20513),
    .in2(net_20514_cascademuxed),
    .in3(gnd),
    .lcout(net_16582),
    .ltout(),
    .sr(net_20530)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_4_17_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_21020),
    .clk(net_21021),
    .in0(gnd),
    .in1(gnd),
    .in2(net_20982_cascademuxed),
    .in3(gnd),
    .lcout(net_17070),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_4_18_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_21097),
    .in1(net_21098),
    .in2(net_21099_cascademuxed),
    .in3(net_21100),
    .lcout(net_17192),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_4_18_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21144),
    .in0(net_21109),
    .in1(gnd),
    .in2(net_21111_cascademuxed),
    .in3(net_21112),
    .lcout(net_17194),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_4_18_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_21133),
    .in1(net_21134),
    .in2(net_21135_cascademuxed),
    .in3(net_21136),
    .lcout(net_17198),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_4_18_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_21144),
    .in0(net_21139),
    .in1(gnd),
    .in2(net_21141_cascademuxed),
    .in3(gnd),
    .lcout(net_17199),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_19_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_21226),
    .in1(net_21227),
    .in2(net_21228_cascademuxed),
    .in3(net_21229),
    .lcout(net_17316),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_19_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_21232),
    .in1(net_21233),
    .in2(net_21234_cascademuxed),
    .in3(net_21235),
    .lcout(net_17317),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_19_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_21244),
    .in1(net_21245),
    .in2(net_21246_cascademuxed),
    .in3(net_21247),
    .lcout(net_17319),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_4_20_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_21349),
    .in1(net_21350),
    .in2(net_21351_cascademuxed),
    .in3(net_21352),
    .lcout(net_17439),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_5_12_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_24236),
    .clk(net_24237),
    .in0(net_24202),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_20287),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_20_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_25220),
    .clk(net_25221),
    .in0(gnd),
    .in1(gnd),
    .in2(net_25188_cascademuxed),
    .in3(gnd),
    .lcout(net_21271),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_5_5_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_23376),
    .in0(gnd),
    .in1(gnd),
    .in2(net_23331_cascademuxed),
    .in3(gnd),
    .lcout(net_19424),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_11_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_0 (
    .carryin(t46),
    .carryout(t48),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_31223_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_1 (
    .carryin(t48),
    .carryout(net_31226),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_31228),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_7_12_2 (
    .carryin(net_31226),
    .carryout(net_31232),
    .ce(),
    .clk(net_31268),
    .in0(gnd),
    .in1(net_31234),
    .in2(gnd),
    .in3(net_31236),
    .lcout(net_27687),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_7_12_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_31268),
    .in0(net_31239),
    .in1(gnd),
    .in2(gnd),
    .in3(net_31242),
    .lcout(net_27688),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_12_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_31251),
    .in1(net_31252),
    .in2(net_31253_cascademuxed),
    .in3(net_31254),
    .lcout(net_27690),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000100010000),
    .SEQ_MODE(4'b0000)
  ) lc40_7_1_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_29836_cascademuxed),
    .in3(net_29837),
    .lcout(net_26554),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_10_0 (
    .carryin(t50),
    .carryout(t52),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34807),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_10_1 (
    .carryin(t52),
    .carryout(net_34811),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34813),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_10_2 (
    .carryin(net_34811),
    .carryout(net_34817),
    .ce(),
    .clk(net_34853),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34820_cascademuxed),
    .in3(net_34821),
    .lcout(net_30903),
    .ltout(),
    .sr(net_34854)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_10_3 (
    .carryin(net_34817),
    .carryout(net_34823),
    .ce(),
    .clk(net_34853),
    .in0(gnd),
    .in1(net_34825),
    .in2(gnd),
    .in3(net_34827),
    .lcout(net_30904),
    .ltout(),
    .sr(net_34854)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_10_4 (
    .carryin(net_34823),
    .carryout(net_34829),
    .ce(),
    .clk(net_34853),
    .in0(gnd),
    .in1(net_34831),
    .in2(gnd),
    .in3(net_34833),
    .lcout(net_30905),
    .ltout(),
    .sr(net_34854)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_10_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_34853),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34838_cascademuxed),
    .in3(net_34839),
    .lcout(net_30906),
    .ltout(),
    .sr(net_34854)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_34842),
    .in1(net_34843),
    .in2(net_34844_cascademuxed),
    .in3(net_34845),
    .lcout(net_30907),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_34849),
    .in2(net_34850_cascademuxed),
    .in3(net_34851),
    .lcout(net_30908),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_8_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_34975),
    .clk(net_34976),
    .in0(gnd),
    .in1(gnd),
    .in2(net_34961_cascademuxed),
    .in3(gnd),
    .lcout(net_31029),
    .ltout(),
    .sr(net_34977)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35099),
    .in0(net_35058),
    .in1(gnd),
    .in2(net_35060_cascademuxed),
    .in3(gnd),
    .lcout(net_31148),
    .ltout(),
    .sr(net_35100)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_8_17_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_35714),
    .in0(gnd),
    .in1(gnd),
    .in2(net_35699_cascademuxed),
    .in3(gnd),
    .lcout(net_31767),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_23_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_36452),
    .in0(net_36435),
    .in1(net_36436),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_32505),
    .ltout(),
    .sr(net_36453)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b1000)
  ) lc40_8_24_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_36574),
    .clk(net_36575),
    .in0(net_36564),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_32629),
    .ltout(),
    .sr(net_36576)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_24_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_25_0 (
    .carryin(t55),
    .carryout(t57),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_36652),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_25_1 (
    .carryin(t57),
    .carryout(net_36656),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_36658),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_25_2 (
    .carryin(net_36656),
    .carryout(net_36662),
    .ce(),
    .clk(net_36698),
    .in0(gnd),
    .in1(gnd),
    .in2(net_36665_cascademuxed),
    .in3(net_36666),
    .lcout(net_32748),
    .ltout(),
    .sr(net_36699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_25_3 (
    .carryin(net_36662),
    .carryout(net_36668),
    .ce(),
    .clk(net_36698),
    .in0(gnd),
    .in1(gnd),
    .in2(net_36671_cascademuxed),
    .in3(net_36672),
    .lcout(net_32749),
    .ltout(),
    .sr(net_36699)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_25_4 (
    .carryin(net_36668),
    .carryout(net_36674),
    .ce(),
    .clk(net_36698),
    .in0(gnd),
    .in1(net_36676),
    .in2(gnd),
    .in3(net_36678),
    .lcout(net_32750),
    .ltout(),
    .sr(net_36699)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b1000)
  ) lc40_8_25_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(net_36698),
    .in0(gnd),
    .in1(net_36682),
    .in2(gnd),
    .in3(net_36684),
    .lcout(net_32751),
    .ltout(),
    .sr(net_36699)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_25_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_36687),
    .in1(net_36688),
    .in2(net_36689_cascademuxed),
    .in3(gnd),
    .lcout(net_32752),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_25_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_36693),
    .in1(net_36694),
    .in2(net_36695_cascademuxed),
    .in3(net_36696),
    .lcout(net_32753),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000001000000011),
    .SEQ_MODE(4'b0000)
  ) lc40_8_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33828),
    .in1(gnd),
    .in2(net_33830_cascademuxed),
    .in3(net_33831),
    .lcout(net_29882),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_33868),
    .clk(net_33869),
    .in0(gnd),
    .in1(net_33835),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_29883),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_8_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33840),
    .in1(net_33841),
    .in2(net_33842_cascademuxed),
    .in3(net_33843),
    .lcout(net_29884),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_33847),
    .in2(net_33848_cascademuxed),
    .in3(net_33849),
    .lcout(net_29885),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011011100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33852),
    .in1(net_33853),
    .in2(net_33854_cascademuxed),
    .in3(net_33855),
    .lcout(net_29886),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110100111010001),
    .SEQ_MODE(4'b0000)
  ) lc40_8_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33858),
    .in1(net_33859),
    .in2(net_33860_cascademuxed),
    .in3(net_33861),
    .lcout(net_29887),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0011011000111100),
    .SEQ_MODE(4'b0000)
  ) lc40_8_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33864),
    .in1(net_33865),
    .in2(net_33866_cascademuxed),
    .in3(net_33867),
    .lcout(net_29888),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_8_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_33952),
    .in2(gnd),
    .in3(net_33954),
    .lcout(net_30041),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1010101010000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33969),
    .in1(net_33970),
    .in2(net_33971_cascademuxed),
    .in3(net_33972),
    .lcout(net_30044),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0010010000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_8_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_33991),
    .clk(net_33992),
    .in0(net_33975),
    .in1(net_33976),
    .in2(net_33977_cascademuxed),
    .in3(net_33978),
    .lcout(net_30045),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110101111111111),
    .SEQ_MODE(4'b0000)
  ) lc40_8_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33981),
    .in1(net_33982),
    .in2(net_33983_cascademuxed),
    .in3(net_33984),
    .lcout(net_30046),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b0000)
  ) lc40_8_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_33987),
    .in1(net_33988),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30047),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_8_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_30164),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_8_9_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_10_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_38643),
    .in1(net_38644),
    .in2(net_38645_cascademuxed),
    .in3(net_38646),
    .lcout(net_34733),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38683),
    .clk(net_38684),
    .in0(net_38649),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34734),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_9_10_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_38661),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34736),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_10_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_38673),
    .in1(net_38674),
    .in2(net_38675_cascademuxed),
    .in3(net_38676),
    .lcout(net_34738),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_10_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38683),
    .clk(net_38684),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38681_cascademuxed),
    .in3(gnd),
    .lcout(net_34739),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_11_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38806),
    .clk(net_38807),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_38793),
    .lcout(net_34860),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_12_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38929),
    .clk(net_38930),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38891_cascademuxed),
    .in3(gnd),
    .lcout(net_34979),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_18_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39667),
    .clk(net_39668),
    .in0(gnd),
    .in1(gnd),
    .in2(net_39629_cascademuxed),
    .in3(gnd),
    .lcout(net_35717),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_18_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_39667),
    .clk(net_39668),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(net_39654),
    .lcout(net_35721),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_27_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_40734),
    .in1(gnd),
    .in2(net_40736_cascademuxed),
    .in3(gnd),
    .lcout(net_36824),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_27_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_40774),
    .clk(net_40775),
    .in0(gnd),
    .in1(gnd),
    .in2(net_40760_cascademuxed),
    .in3(net_40761),
    .lcout(net_36828),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b1000)
  ) lc40_9_27_7 (
    .carryin(gnd),
    .carryout(),
    .ce(net_40774),
    .clk(net_40775),
    .in0(net_40770),
    .in1(net_40771),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_36830),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_28_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_40857),
    .in1(gnd),
    .in2(net_40859_cascademuxed),
    .in3(gnd),
    .lcout(net_36947),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_28_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_40864),
    .in2(net_40865_cascademuxed),
    .in3(net_40866),
    .lcout(net_36948),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_9_28_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_40882),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_36951),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1001010110001101),
    .SEQ_MODE(4'b1000)
  ) lc40_9_28_6 (
    .carryin(gnd),
    .carryout(),
    .ce(net_40897),
    .clk(net_40898),
    .in0(net_40887),
    .in1(net_40888),
    .in2(net_40889_cascademuxed),
    .in3(net_40890),
    .lcout(net_36952),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110110111111111),
    .SEQ_MODE(4'b0000)
  ) lc40_9_29_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_40974),
    .in1(net_40975),
    .in2(net_40976_cascademuxed),
    .in3(net_40977),
    .lcout(net_37069),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000100000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_29_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_40993),
    .in2(gnd),
    .in3(net_40995),
    .lcout(net_37072),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b0000)
  ) lc40_9_29_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_41004),
    .in1(net_41005),
    .in2(net_41006_cascademuxed),
    .in3(net_41007),
    .lcout(net_37074),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1100001001110011),
    .SEQ_MODE(4'b1000)
  ) lc40_9_2_0 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37699),
    .clk(net_37700),
    .in0(net_37653),
    .in1(net_37654),
    .in2(net_37655_cascademuxed),
    .in3(net_37656),
    .lcout(net_33712),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_2_1 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37659),
    .in1(gnd),
    .in2(net_37661_cascademuxed),
    .in3(net_37662),
    .lcout(net_33713),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_2_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37665),
    .in1(net_37666),
    .in2(net_37667_cascademuxed),
    .in3(net_37668),
    .lcout(net_33714),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_2_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_37673_cascademuxed),
    .in3(net_37674),
    .lcout(net_33715),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_2_4 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37677),
    .in1(net_37678),
    .in2(net_37679_cascademuxed),
    .in3(net_37680),
    .lcout(net_33716),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_9_2_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_37684),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_33717),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001001100110011),
    .SEQ_MODE(4'b0000)
  ) lc40_9_2_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37689),
    .in1(net_37690),
    .in2(net_37691_cascademuxed),
    .in3(net_37692),
    .lcout(net_33718),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000010000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_2_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_37696),
    .in2(gnd),
    .in3(net_37698),
    .lcout(net_33719),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1110100011010011),
    .SEQ_MODE(4'b0000)
  ) lc40_9_30_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_41097),
    .in1(net_41098),
    .in2(net_41099_cascademuxed),
    .in3(net_41100),
    .lcout(net_37192),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101010101101010),
    .SEQ_MODE(4'b0000)
  ) lc40_9_30_2 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_41109),
    .in1(net_41110),
    .in2(net_41111_cascademuxed),
    .in3(net_41112),
    .lcout(net_37194),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_30_5 (
    .carryin(gnd),
    .carryout(),
    .ce(net_41143),
    .clk(net_41144),
    .in0(net_41127),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_37197),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000111000001100),
    .SEQ_MODE(4'b0000)
  ) lc40_9_30_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_41139),
    .in1(net_41140),
    .in2(gnd),
    .in3(net_41142),
    .lcout(net_37199),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000001000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_3_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37776),
    .in1(net_37777),
    .in2(net_37778_cascademuxed),
    .in3(net_37779),
    .lcout(net_33871),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0101000100010001),
    .SEQ_MODE(4'b1000)
  ) lc40_9_3_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37822),
    .clk(net_37823),
    .in0(gnd),
    .in1(net_37783),
    .in2(net_37784_cascademuxed),
    .in3(net_37785),
    .lcout(net_33872),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000001101100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_3_2 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37822),
    .clk(net_37823),
    .in0(net_37788),
    .in1(net_37789),
    .in2(net_37790_cascademuxed),
    .in3(net_37791),
    .lcout(net_33873),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000001),
    .SEQ_MODE(4'b0000)
  ) lc40_9_3_3 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37794),
    .in1(net_37795),
    .in2(net_37796_cascademuxed),
    .in3(net_37797),
    .lcout(net_33874),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b1111111111111101),
    .SEQ_MODE(4'b1000)
  ) lc40_9_3_4 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37822),
    .clk(net_37823),
    .in0(net_37800),
    .in1(net_37801),
    .in2(net_37802_cascademuxed),
    .in3(net_37803),
    .lcout(net_33875),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0001000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_3_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37806),
    .in1(net_37807),
    .in2(net_37808_cascademuxed),
    .in3(net_37809),
    .lcout(net_33876),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000101000101),
    .SEQ_MODE(4'b0000)
  ) lc40_9_3_6 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37812),
    .in1(net_37813),
    .in2(net_37814_cascademuxed),
    .in3(net_37815),
    .lcout(net_33877),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000010000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_3_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37818),
    .in1(net_37819),
    .in2(net_37820_cascademuxed),
    .in3(net_37821),
    .lcout(net_33878),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_4_0 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37899),
    .in1(gnd),
    .in2(net_37901_cascademuxed),
    .in3(gnd),
    .lcout(net_33994),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000010),
    .SEQ_MODE(4'b1000)
  ) lc40_9_4_1 (
    .carryin(gnd),
    .carryout(),
    .ce(net_37945),
    .clk(net_37946),
    .in0(net_37905),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_33995),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000100011),
    .SEQ_MODE(4'b0000)
  ) lc40_9_4_5 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(net_37929),
    .in1(net_37930),
    .in2(net_37931_cascademuxed),
    .in3(gnd),
    .lcout(net_33999),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000100),
    .SEQ_MODE(4'b1000)
  ) lc40_9_5_3 (
    .carryin(gnd),
    .carryout(),
    .ce(net_38068),
    .clk(net_38069),
    .in0(gnd),
    .in1(net_38041),
    .in2(gnd),
    .in3(gnd),
    .lcout(net_34120),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_7_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_0 (
    .carryin(t67),
    .carryout(t69),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38393_cascademuxed),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0000000000000000),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_1 (
    .carryin(t69),
    .carryout(net_38396),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_38398),
    .in2(gnd),
    .in3(gnd),
    .lcout(),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_2 (
    .carryin(net_38396),
    .carryout(net_38402),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38405_cascademuxed),
    .in3(net_38406),
    .lcout(net_34488),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_3 (
    .carryin(net_38402),
    .carryout(net_38408),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38411_cascademuxed),
    .in3(net_38412),
    .lcout(net_34489),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_4 (
    .carryin(net_38408),
    .carryout(net_38414),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38417_cascademuxed),
    .in3(net_38418),
    .lcout(net_34490),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_5 (
    .carryin(net_38414),
    .carryout(net_38420),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38423_cascademuxed),
    .in3(net_38424),
    .lcout(net_34491),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b1),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_6 (
    .carryin(net_38420),
    .carryout(net_38426),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(gnd),
    .in2(net_38429_cascademuxed),
    .in3(net_38430),
    .lcout(net_34492),
    .ltout(),
    .sr(gnd)
  );
  LogicCell40 #(
    .C_ON(1'b0),
    .LUT_INIT(16'b0110100110010110),
    .SEQ_MODE(4'b0000)
  ) lc40_9_8_7 (
    .carryin(gnd),
    .carryout(),
    .ce(),
    .clk(gnd),
    .in0(gnd),
    .in1(net_38434),
    .in2(gnd),
    .in3(net_38436),
    .lcout(net_34493),
    .ltout(),
    .sr(gnd)
  );
  Odrv4 odrv_10_10_38565_31037 (
    .I(net_38565),
    .O(net_31037)
  );
  Odrv4 odrv_10_10_38565_42535 (
    .I(net_38565),
    .O(net_42535)
  );
  Odrv4 odrv_10_11_38688_42665 (
    .I(net_38688),
    .O(net_42665)
  );
  Odrv4 odrv_10_12_38811_42781 (
    .I(net_38811),
    .O(net_42781)
  );
  Odrv4 odrv_10_12_38812_42783 (
    .I(net_38812),
    .O(net_42783)
  );
  Odrv4 odrv_10_12_38813_42785 (
    .I(net_38813),
    .O(net_42785)
  );
  Odrv4 odrv_10_12_38815_38945 (
    .I(net_38815),
    .O(net_38945)
  );
  Odrv4 odrv_10_13_38932_42898 (
    .I(net_38932),
    .O(net_42898)
  );
  Odrv4 odrv_10_13_38935_42906 (
    .I(net_38935),
    .O(net_42906)
  );
  Odrv4 odrv_10_14_39057_43027 (
    .I(net_39057),
    .O(net_43027)
  );
  Odrv4 odrv_10_14_39060_42674 (
    .I(net_39060),
    .O(net_42674)
  );
  Odrv4 odrv_10_15_39178_38957 (
    .I(net_39178),
    .O(net_38957)
  );
  Odrv4 odrv_10_15_39180_43150 (
    .I(net_39180),
    .O(net_43150)
  );
  Odrv4 odrv_10_15_39182_38965 (
    .I(net_39182),
    .O(net_38965)
  );
  Odrv4 odrv_10_17_39426_39207 (
    .I(net_39426),
    .O(net_39207)
  );
  Odrv4 odrv_10_17_39426_39570 (
    .I(net_39426),
    .O(net_39570)
  );
  Odrv4 odrv_10_17_39426_43037 (
    .I(net_39426),
    .O(net_43037)
  );
  Odrv4 odrv_10_17_39426_43403 (
    .I(net_39426),
    .O(net_43403)
  );
  Odrv4 odrv_10_17_39427_39209 (
    .I(net_39427),
    .O(net_39209)
  );
  Odrv4 odrv_10_17_39427_43398 (
    .I(net_39427),
    .O(net_43398)
  );
  Odrv4 odrv_10_17_39427_43405 (
    .I(net_39427),
    .O(net_43405)
  );
  Odrv4 odrv_10_17_39428_39211 (
    .I(net_39428),
    .O(net_39211)
  );
  Odrv4 odrv_10_17_39428_43041 (
    .I(net_39428),
    .O(net_43041)
  );
  Odrv4 odrv_10_17_39428_43279 (
    .I(net_39428),
    .O(net_43279)
  );
  Odrv4 odrv_10_17_39428_43400 (
    .I(net_39428),
    .O(net_43400)
  );
  Odrv4 odrv_10_17_39428_43407 (
    .I(net_39428),
    .O(net_43407)
  );
  Odrv4 odrv_10_17_39429_35732 (
    .I(net_39429),
    .O(net_35732)
  );
  Odrv4 odrv_10_17_39429_39213 (
    .I(net_39429),
    .O(net_39213)
  );
  Odrv4 odrv_10_17_39429_39577 (
    .I(net_39429),
    .O(net_39577)
  );
  Odrv4 odrv_10_17_39429_43043 (
    .I(net_39429),
    .O(net_43043)
  );
  Odrv4 odrv_10_17_39429_43281 (
    .I(net_39429),
    .O(net_43281)
  );
  Odrv4 odrv_10_17_39430_35734 (
    .I(net_39430),
    .O(net_35734)
  );
  Odrv4 odrv_10_17_39430_39325 (
    .I(net_39430),
    .O(net_39325)
  );
  Odrv4 odrv_10_17_39430_39579 (
    .I(net_39430),
    .O(net_39579)
  );
  Odrv4 odrv_10_17_39430_43157 (
    .I(net_39430),
    .O(net_43157)
  );
  Odrv4 odrv_10_17_39430_43283 (
    .I(net_39430),
    .O(net_43283)
  );
  Odrv4 odrv_10_17_39431_39327 (
    .I(net_39431),
    .O(net_39327)
  );
  Odrv4 odrv_10_17_39431_39455 (
    .I(net_39431),
    .O(net_39455)
  );
  Odrv4 odrv_10_17_39431_39564 (
    .I(net_39431),
    .O(net_39564)
  );
  Odrv4 odrv_10_17_39431_43159 (
    .I(net_39431),
    .O(net_43159)
  );
  Odrv4 odrv_10_17_39431_43285 (
    .I(net_39431),
    .O(net_43285)
  );
  Odrv4 odrv_10_18_39547_35861 (
    .I(net_39547),
    .O(net_35861)
  );
  Odrv4 odrv_10_18_39547_39326 (
    .I(net_39547),
    .O(net_39326)
  );
  Odrv4 odrv_10_18_39547_39689 (
    .I(net_39547),
    .O(net_39689)
  );
  Odrv4 odrv_10_18_39547_43156 (
    .I(net_39547),
    .O(net_43156)
  );
  Odrv4 odrv_10_18_39548_35853 (
    .I(net_39548),
    .O(net_35853)
  );
  Odrv4 odrv_10_18_39548_39328 (
    .I(net_39548),
    .O(net_39328)
  );
  Odrv4 odrv_10_18_39548_39691 (
    .I(net_39548),
    .O(net_39691)
  );
  Odrv4 odrv_10_18_39548_43158 (
    .I(net_39548),
    .O(net_43158)
  );
  Odrv4 odrv_10_18_39548_43286 (
    .I(net_39548),
    .O(net_43286)
  );
  Odrv4 odrv_10_18_39549_39330 (
    .I(net_39549),
    .O(net_39330)
  );
  Odrv4 odrv_10_18_39549_43160 (
    .I(net_39549),
    .O(net_43160)
  );
  Odrv4 odrv_10_18_39549_43519 (
    .I(net_39549),
    .O(net_43519)
  );
  Odrv4 odrv_10_18_39549_43526 (
    .I(net_39549),
    .O(net_43526)
  );
  Odrv4 odrv_10_18_39550_39332 (
    .I(net_39550),
    .O(net_39332)
  );
  Odrv4 odrv_10_18_39550_39685 (
    .I(net_39550),
    .O(net_39685)
  );
  Odrv4 odrv_10_18_39550_43290 (
    .I(net_39550),
    .O(net_43290)
  );
  Odrv4 odrv_10_18_39550_43528 (
    .I(net_39550),
    .O(net_43528)
  );
  Odrv4 odrv_10_18_39551_35851 (
    .I(net_39551),
    .O(net_35851)
  );
  Odrv4 odrv_10_18_39551_39334 (
    .I(net_39551),
    .O(net_39334)
  );
  Odrv4 odrv_10_18_39551_43164 (
    .I(net_39551),
    .O(net_43164)
  );
  Odrv4 odrv_10_18_39551_43523 (
    .I(net_39551),
    .O(net_43523)
  );
  Odrv4 odrv_10_18_39552_35855 (
    .I(net_39552),
    .O(net_35855)
  );
  Odrv4 odrv_10_18_39552_39336 (
    .I(net_39552),
    .O(net_39336)
  );
  Odrv4 odrv_10_18_39552_43166 (
    .I(net_39552),
    .O(net_43166)
  );
  Odrv4 odrv_10_18_39552_43532 (
    .I(net_39552),
    .O(net_43532)
  );
  Odrv4 odrv_10_18_39553_39448 (
    .I(net_39553),
    .O(net_39448)
  );
  Odrv4 odrv_10_18_39553_43280 (
    .I(net_39553),
    .O(net_43280)
  );
  Odrv4 odrv_10_18_39553_43534 (
    .I(net_39553),
    .O(net_43534)
  );
  Odrv4 odrv_10_18_39554_39687 (
    .I(net_39554),
    .O(net_39687)
  );
  Odrv4 odrv_10_18_39554_43282 (
    .I(net_39554),
    .O(net_43282)
  );
  Odrv4 odrv_10_18_39554_43408 (
    .I(net_39554),
    .O(net_43408)
  );
  Odrv4 odrv_10_19_39670_39812 (
    .I(net_39670),
    .O(net_39812)
  );
  Odrv4 odrv_10_19_39670_43636 (
    .I(net_39670),
    .O(net_43636)
  );
  Odrv4 odrv_10_19_39671_35976 (
    .I(net_39671),
    .O(net_35976)
  );
  Odrv4 odrv_10_19_39671_43640 (
    .I(net_39671),
    .O(net_43640)
  );
  Odrv4 odrv_10_19_39672_39816 (
    .I(net_39672),
    .O(net_39816)
  );
  Odrv4 odrv_10_19_39672_43411 (
    .I(net_39672),
    .O(net_43411)
  );
  Odrv4 odrv_10_19_39672_43642 (
    .I(net_39672),
    .O(net_43642)
  );
  Odrv4 odrv_10_19_39673_43413 (
    .I(net_39673),
    .O(net_43413)
  );
  Odrv4 odrv_10_19_39673_43644 (
    .I(net_39673),
    .O(net_43644)
  );
  Odrv4 odrv_10_19_39674_35974 (
    .I(net_39674),
    .O(net_35974)
  );
  Odrv4 odrv_10_19_39674_43646 (
    .I(net_39674),
    .O(net_43646)
  );
  Odrv4 odrv_10_19_39675_43638 (
    .I(net_39675),
    .O(net_43638)
  );
  Odrv4 odrv_10_19_39676_35980 (
    .I(net_39676),
    .O(net_35980)
  );
  Odrv4 odrv_10_19_39676_39806 (
    .I(net_39676),
    .O(net_39806)
  );
  Odrv4 odrv_10_19_39677_39810 (
    .I(net_39677),
    .O(net_39810)
  );
  Odrv4 odrv_10_20_39793_43759 (
    .I(net_39793),
    .O(net_43759)
  );
  Odrv4 odrv_10_20_39794_43763 (
    .I(net_39794),
    .O(net_43763)
  );
  Odrv12 odrv_10_20_39795_21400 (
    .I(net_39795),
    .O(net_21400)
  );
  Odrv4 odrv_10_20_39795_43765 (
    .I(net_39795),
    .O(net_43765)
  );
  Odrv4 odrv_10_20_39796_39931 (
    .I(net_39796),
    .O(net_39931)
  );
  Odrv4 odrv_10_20_39796_43767 (
    .I(net_39796),
    .O(net_43767)
  );
  Odrv12 odrv_10_26_40533_44250 (
    .I(net_40533),
    .O(net_44250)
  );
  Odrv4 odrv_10_28_40782_40804 (
    .I(net_40782),
    .O(net_40804)
  );
  Odrv4 odrv_10_29_40906_40801 (
    .I(net_40906),
    .O(net_40801)
  );
  Odrv4 odrv_10_7_38199_37983 (
    .I(net_38199),
    .O(net_37983)
  );
  Odrv4 odrv_10_7_38199_41813 (
    .I(net_38199),
    .O(net_41813)
  );
  Odrv4 odrv_10_7_38199_42051 (
    .I(net_38199),
    .O(net_42051)
  );
  Odrv4 odrv_10_7_38199_42162 (
    .I(net_38199),
    .O(net_42162)
  );
  Odrv4 odrv_10_8_38318_42182 (
    .I(net_38318),
    .O(net_42182)
  );
  Odrv4 odrv_11_10_42394_46257 (
    .I(net_42394),
    .O(net_46257)
  );
  Odrv4 odrv_11_10_42397_46375 (
    .I(net_42397),
    .O(net_46375)
  );
  Odrv4 odrv_11_10_42398_38698 (
    .I(net_42398),
    .O(net_38698)
  );
  Odrv4 odrv_11_10_42398_42419 (
    .I(net_42398),
    .O(net_42419)
  );
  Odrv4 odrv_11_10_42398_42545 (
    .I(net_42398),
    .O(net_42545)
  );
  Odrv4 odrv_11_10_42398_46011 (
    .I(net_42398),
    .O(net_46011)
  );
  Odrv4 odrv_11_10_42398_46249 (
    .I(net_42398),
    .O(net_46249)
  );
  Odrv4 odrv_11_10_42398_46370 (
    .I(net_42398),
    .O(net_46370)
  );
  Odrv4 odrv_11_10_42398_46377 (
    .I(net_42398),
    .O(net_46377)
  );
  Odrv4 odrv_11_10_42400_42295 (
    .I(net_42400),
    .O(net_42295)
  );
  Odrv4 odrv_11_10_42400_42530 (
    .I(net_42400),
    .O(net_42530)
  );
  Odrv4 odrv_11_10_42400_42549 (
    .I(net_42400),
    .O(net_42549)
  );
  Odrv4 odrv_11_10_42400_46127 (
    .I(net_42400),
    .O(net_46127)
  );
  Odrv4 odrv_11_10_42400_46253 (
    .I(net_42400),
    .O(net_46253)
  );
  Odrv4 odrv_11_10_42401_42534 (
    .I(net_42401),
    .O(net_42534)
  );
  Odrv4 odrv_11_10_42401_46255 (
    .I(net_42401),
    .O(net_46255)
  );
  Odrv4 odrv_11_10_42401_46383 (
    .I(net_42401),
    .O(net_46383)
  );
  Odrv4 odrv_11_12_42641_46610 (
    .I(net_42641),
    .O(net_46610)
  );
  Odrv4 odrv_11_12_42642_42786 (
    .I(net_42642),
    .O(net_42786)
  );
  Odrv4 odrv_11_12_42643_46614 (
    .I(net_42643),
    .O(net_46614)
  );
  Odrv4 odrv_11_12_42644_46616 (
    .I(net_42644),
    .O(net_46616)
  );
  Odrv4 odrv_11_12_42647_42780 (
    .I(net_42647),
    .O(net_42780)
  );
  Odrv4 odrv_11_13_42763_39077 (
    .I(net_42763),
    .O(net_39077)
  );
  Odrv4 odrv_11_13_42764_46733 (
    .I(net_42764),
    .O(net_46733)
  );
  Odrv4 odrv_11_13_42765_46735 (
    .I(net_42765),
    .O(net_46735)
  );
  Odrv4 odrv_11_13_42767_39067 (
    .I(net_42767),
    .O(net_39067)
  );
  Odrv12 odrv_11_13_42768_42895 (
    .I(net_42768),
    .O(net_42895)
  );
  Odrv4 odrv_11_13_42769_42899 (
    .I(net_42769),
    .O(net_42899)
  );
  Odrv4 odrv_11_14_42887_46856 (
    .I(net_42887),
    .O(net_46856)
  );
  Odrv4 odrv_11_14_42891_46743 (
    .I(net_42891),
    .O(net_46743)
  );
  Odrv4 odrv_11_14_42893_43026 (
    .I(net_42893),
    .O(net_43026)
  );
  Odrv4 odrv_11_15_43012_42794 (
    .I(net_43012),
    .O(net_42794)
  );
  Odrv4 odrv_11_16_43137_46751 (
    .I(net_43137),
    .O(net_46751)
  );
  Odrv4 odrv_11_16_43137_47100 (
    .I(net_43137),
    .O(net_47100)
  );
  Odrv4 odrv_11_16_43137_47117 (
    .I(net_43137),
    .O(net_47117)
  );
  Odrv4 odrv_11_17_43256_43162 (
    .I(net_43256),
    .O(net_43162)
  );
  Odrv4 odrv_11_17_43256_43399 (
    .I(net_43256),
    .O(net_43399)
  );
  Odrv4 odrv_11_17_43256_47120 (
    .I(net_43256),
    .O(net_47120)
  );
  Odrv4 odrv_11_17_43256_47225 (
    .I(net_43256),
    .O(net_47225)
  );
  Odrv4 odrv_11_18_43379_47348 (
    .I(net_43379),
    .O(net_47348)
  );
  Odrv4 odrv_11_18_43380_47350 (
    .I(net_43380),
    .O(net_47350)
  );
  Odrv4 odrv_11_19_43504_47475 (
    .I(net_43504),
    .O(net_47475)
  );
  Odrv4 odrv_11_20_43626_47596 (
    .I(net_43626),
    .O(net_47596)
  );
  Odrv4 odrv_11_20_43630_43760 (
    .I(net_43630),
    .O(net_43760)
  );
  Odrv4 odrv_11_23_43999_44148 (
    .I(net_43999),
    .O(net_44148)
  );
  Odrv4 odrv_11_23_43999_47726 (
    .I(net_43999),
    .O(net_47726)
  );
  Odrv4 odrv_11_29_44736_44520 (
    .I(net_44736),
    .O(net_44520)
  );
  Odrv4 odrv_11_30_44855_41156 (
    .I(net_44855),
    .O(net_41156)
  );
  Odrv4 odrv_11_30_44857_48824 (
    .I(net_44857),
    .O(net_48824)
  );
  Odrv4 odrv_11_7_42025_45762 (
    .I(net_42025),
    .O(net_45762)
  );
  Odrv4 odrv_11_9_42271_42413 (
    .I(net_42271),
    .O(net_42413)
  );
  Odrv4 odrv_11_9_42272_38577 (
    .I(net_42272),
    .O(net_38577)
  );
  Odrv4 odrv_11_9_42274_42409 (
    .I(net_42274),
    .O(net_42409)
  );
  Odrv4 odrv_12_11_46349_50318 (
    .I(net_46349),
    .O(net_50318)
  );
  Odrv4 odrv_12_11_46351_50091 (
    .I(net_46351),
    .O(net_50091)
  );
  Odrv4 odrv_12_12_46473_50443 (
    .I(net_46473),
    .O(net_50443)
  );
  Odrv4 odrv_12_14_46719_50689 (
    .I(net_46719),
    .O(net_50689)
  );
  Odrv4 odrv_12_14_46721_46504 (
    .I(net_46721),
    .O(net_46504)
  );
  Odrv4 odrv_12_14_46724_46857 (
    .I(net_46724),
    .O(net_46857)
  );
  Odrv4 odrv_12_15_46841_50451 (
    .I(net_46841),
    .O(net_50451)
  );
  Odrv4 odrv_12_15_46842_50812 (
    .I(net_46842),
    .O(net_50812)
  );
  Odrv4 odrv_12_15_46843_46625 (
    .I(net_46843),
    .O(net_46625)
  );
  Odrv4 odrv_12_15_46847_43152 (
    .I(net_46847),
    .O(net_43152)
  );
  Odrv4 odrv_12_16_46967_50939 (
    .I(net_46967),
    .O(net_50939)
  );
  Odrv4 odrv_12_17_47091_51054 (
    .I(net_47091),
    .O(net_51054)
  );
  Odrv4 odrv_12_18_47209_47351 (
    .I(net_47209),
    .O(net_47351)
  );
  Odrv4 odrv_12_18_47209_51175 (
    .I(net_47209),
    .O(net_51175)
  );
  Odrv4 odrv_12_19_47334_51304 (
    .I(net_47334),
    .O(net_51304)
  );
  Odrv4 odrv_12_19_47334_51311 (
    .I(net_47334),
    .O(net_51311)
  );
  Odrv4 odrv_12_21_47578_43892 (
    .I(net_47578),
    .O(net_43892)
  );
  Odrv4 odrv_12_21_47578_47357 (
    .I(net_47578),
    .O(net_47357)
  );
  Odrv4 odrv_12_21_47578_47483 (
    .I(net_47578),
    .O(net_47483)
  );
  Odrv4 odrv_12_21_47578_47720 (
    .I(net_47578),
    .O(net_47720)
  );
  Odrv4 odrv_12_21_47578_51187 (
    .I(net_47578),
    .O(net_51187)
  );
  Odrv4 odrv_12_21_47578_51315 (
    .I(net_47578),
    .O(net_51315)
  );
  Odrv4 odrv_12_21_47578_51544 (
    .I(net_47578),
    .O(net_51544)
  );
  Odrv4 odrv_12_21_47580_47361 (
    .I(net_47580),
    .O(net_47361)
  );
  Odrv4 odrv_12_21_47580_47724 (
    .I(net_47580),
    .O(net_47724)
  );
  Odrv12 odrv_12_21_47580_50313 (
    .I(net_47580),
    .O(net_50313)
  );
  Odrv4 odrv_12_21_47580_51191 (
    .I(net_47580),
    .O(net_51191)
  );
  Odrv4 odrv_12_21_47580_51319 (
    .I(net_47580),
    .O(net_51319)
  );
  Odrv4 odrv_12_21_47580_51550 (
    .I(net_47580),
    .O(net_51550)
  );
  Odrv4 odrv_12_21_47582_47365 (
    .I(net_47582),
    .O(net_47365)
  );
  Odrv4 odrv_12_21_47582_51195 (
    .I(net_47582),
    .O(net_51195)
  );
  Odrv4 odrv_12_21_47585_47718 (
    .I(net_47585),
    .O(net_47718)
  );
  Odrv4 odrv_12_23_47824_44138 (
    .I(net_47824),
    .O(net_44138)
  );
  Odrv4 odrv_12_23_47824_47603 (
    .I(net_47824),
    .O(net_47603)
  );
  Odrv4 odrv_12_23_47824_51433 (
    .I(net_47824),
    .O(net_51433)
  );
  Odrv4 odrv_12_27_48322_48452 (
    .I(net_48322),
    .O(net_48452)
  );
  Odrv4 odrv_12_27_48323_48456 (
    .I(net_48323),
    .O(net_48456)
  );
  Odrv4 odrv_12_28_48440_48583 (
    .I(net_48440),
    .O(net_48583)
  );
  Odrv4 odrv_12_30_48691_48817 (
    .I(net_48691),
    .O(net_48817)
  );
  Odrv12 odrv_12_31_48810_51543 (
    .I(net_48810),
    .O(net_51543)
  );
  Odrv4 odrv_12_31_48810_52679 (
    .I(net_48810),
    .O(net_52679)
  );
  Odrv4 odrv_12_8_45980_49949 (
    .I(net_45980),
    .O(net_49949)
  );
  Odrv4 odrv_12_8_45985_38463 (
    .I(net_45985),
    .O(net_38463)
  );
  Odrv4 odrv_13_12_50302_54268 (
    .I(net_50302),
    .O(net_54268)
  );
  Odrv4 odrv_13_12_50305_54276 (
    .I(net_50305),
    .O(net_54276)
  );
  Odrv4 odrv_13_12_50308_46612 (
    .I(net_50308),
    .O(net_46612)
  );
  Odrv4 odrv_13_12_50309_42778 (
    .I(net_50309),
    .O(net_42778)
  );
  Odrv4 odrv_13_13_50425_50567 (
    .I(net_50425),
    .O(net_50567)
  );
  Odrv4 odrv_13_13_50425_54162 (
    .I(net_50425),
    .O(net_54162)
  );
  Odrv4 odrv_13_13_50426_54395 (
    .I(net_50426),
    .O(net_54395)
  );
  Odrv4 odrv_13_13_50427_54397 (
    .I(net_50427),
    .O(net_54397)
  );
  Odrv4 odrv_13_13_50431_42909 (
    .I(net_50431),
    .O(net_42909)
  );
  Odrv4 odrv_13_13_50432_46737 (
    .I(net_50432),
    .O(net_46737)
  );
  Odrv4 odrv_13_14_50548_54514 (
    .I(net_50548),
    .O(net_54514)
  );
  Odrv4 odrv_13_14_50549_54159 (
    .I(net_50549),
    .O(net_54159)
  );
  Odrv4 odrv_13_14_50554_54281 (
    .I(net_50554),
    .O(net_54281)
  );
  Odrv4 odrv_13_15_50671_50813 (
    .I(net_50671),
    .O(net_50813)
  );
  Odrv4 odrv_13_15_50671_54637 (
    .I(net_50671),
    .O(net_54637)
  );
  Odrv4 odrv_13_15_50672_54641 (
    .I(net_50672),
    .O(net_54641)
  );
  Odrv4 odrv_13_15_50674_54414 (
    .I(net_50674),
    .O(net_54414)
  );
  Odrv4 odrv_13_15_50676_46979 (
    .I(net_50676),
    .O(net_46979)
  );
  Odrv4 odrv_13_15_50678_50811 (
    .I(net_50678),
    .O(net_50811)
  );
  Odrv4 odrv_13_16_50796_54407 (
    .I(net_50796),
    .O(net_54407)
  );
  Odrv4 odrv_13_16_50797_54409 (
    .I(net_50797),
    .O(net_54409)
  );
  Odrv4 odrv_13_16_50798_54777 (
    .I(net_50798),
    .O(net_54777)
  );
  Odrv4 odrv_13_16_50799_47102 (
    .I(net_50799),
    .O(net_47102)
  );
  Odrv4 odrv_13_16_50800_54527 (
    .I(net_50800),
    .O(net_54527)
  );
  Odrv4 odrv_13_16_50801_50697 (
    .I(net_50801),
    .O(net_50697)
  );
  Odrv4 odrv_13_17_50917_51059 (
    .I(net_50917),
    .O(net_51059)
  );
  Odrv4 odrv_13_17_50918_50698 (
    .I(net_50918),
    .O(net_50698)
  );
  Odrv4 odrv_13_17_50919_51063 (
    .I(net_50919),
    .O(net_51063)
  );
  Odrv4 odrv_13_17_50920_51055 (
    .I(net_50920),
    .O(net_51055)
  );
  Odrv4 odrv_13_17_50921_54900 (
    .I(net_50921),
    .O(net_54900)
  );
  Odrv4 odrv_13_17_50922_54536 (
    .I(net_50922),
    .O(net_54536)
  );
  Odrv4 odrv_13_17_50924_54652 (
    .I(net_50924),
    .O(net_54652)
  );
  Odrv4 odrv_13_19_51164_51307 (
    .I(net_51164),
    .O(net_51307)
  );
  Odrv4 odrv_13_19_51164_55133 (
    .I(net_51164),
    .O(net_55133)
  );
  Odrv4 odrv_13_19_51167_55018 (
    .I(net_51167),
    .O(net_55018)
  );
  Odrv4 odrv_13_19_51167_55139 (
    .I(net_51167),
    .O(net_55139)
  );
  Odrv4 odrv_13_20_51289_51071 (
    .I(net_51289),
    .O(net_51071)
  );
  Odrv4 odrv_13_21_51415_51310 (
    .I(net_51415),
    .O(net_51310)
  );
  Odrv4 odrv_13_22_51535_51681 (
    .I(net_51535),
    .O(net_51681)
  );
  Odrv4 odrv_13_27_52153_55880 (
    .I(net_52153),
    .O(net_55880)
  );
  Odrv12 odrv_13_31_52639_55128 (
    .I(net_52639),
    .O(net_55128)
  );
  Odrv12 odrv_13_31_52640_55250 (
    .I(net_52640),
    .O(net_55250)
  );
  Odrv4 odrv_13_3_49196_52929 (
    .I(net_49196),
    .O(net_52929)
  );
  Odrv4 odrv_13_8_49816_49946 (
    .I(net_49816),
    .O(net_49946)
  );
  Odrv4 odrv_13_9_49935_53674 (
    .I(net_49935),
    .O(net_53674)
  );
  Odrv4 odrv_14_10_53894_46363 (
    .I(net_53894),
    .O(net_46363)
  );
  Odrv4 odrv_14_11_54012_57981 (
    .I(net_54012),
    .O(net_57981)
  );
  Odrv4 odrv_14_11_54012_57988 (
    .I(net_54012),
    .O(net_57988)
  );
  Odrv4 odrv_14_11_54014_54161 (
    .I(net_54014),
    .O(net_54161)
  );
  Odrv4 odrv_14_12_54133_57995 (
    .I(net_54133),
    .O(net_57995)
  );
  Odrv4 odrv_14_12_54134_58102 (
    .I(net_54134),
    .O(net_58102)
  );
  Odrv4 odrv_14_12_54137_46613 (
    .I(net_54137),
    .O(net_46613)
  );
  Odrv4 odrv_14_12_54138_46615 (
    .I(net_54138),
    .O(net_46615)
  );
  Odrv4 odrv_14_12_54140_57867 (
    .I(net_54140),
    .O(net_57867)
  );
  Odrv4 odrv_14_12_54140_57993 (
    .I(net_54140),
    .O(net_57993)
  );
  Odrv4 odrv_14_13_54256_50570 (
    .I(net_54256),
    .O(net_50570)
  );
  Odrv4 odrv_14_13_54257_58225 (
    .I(net_54257),
    .O(net_58225)
  );
  Odrv4 odrv_14_13_54259_58229 (
    .I(net_54259),
    .O(net_58229)
  );
  Odrv4 odrv_14_13_54259_58236 (
    .I(net_54259),
    .O(net_58236)
  );
  Odrv4 odrv_14_13_54260_50560 (
    .I(net_54260),
    .O(net_50560)
  );
  Odrv4 odrv_14_13_54260_58231 (
    .I(net_54260),
    .O(net_58231)
  );
  Odrv4 odrv_14_13_54261_50564 (
    .I(net_54261),
    .O(net_50564)
  );
  Odrv4 odrv_14_13_54261_58223 (
    .I(net_54261),
    .O(net_58223)
  );
  Odrv4 odrv_14_13_54262_54157 (
    .I(net_54262),
    .O(net_54157)
  );
  Odrv4 odrv_14_13_54263_50568 (
    .I(net_54263),
    .O(net_50568)
  );
  Odrv4 odrv_14_14_54379_58241 (
    .I(net_54379),
    .O(net_58241)
  );
  Odrv4 odrv_14_14_54379_58344 (
    .I(net_54379),
    .O(net_58344)
  );
  Odrv4 odrv_14_14_54381_54288 (
    .I(net_54381),
    .O(net_54288)
  );
  Odrv4 odrv_14_14_54381_54525 (
    .I(net_54381),
    .O(net_54525)
  );
  Odrv4 odrv_14_14_54382_58121 (
    .I(net_54382),
    .O(net_58121)
  );
  Odrv4 odrv_14_14_54383_54166 (
    .I(net_54383),
    .O(net_54166)
  );
  Odrv4 odrv_14_14_54386_54282 (
    .I(net_54386),
    .O(net_54282)
  );
  Odrv4 odrv_14_14_54386_54519 (
    .I(net_54386),
    .O(net_54519)
  );
  Odrv4 odrv_14_15_54503_54283 (
    .I(net_54503),
    .O(net_54283)
  );
  Odrv4 odrv_14_15_54504_54285 (
    .I(net_54504),
    .O(net_54285)
  );
  Odrv4 odrv_14_15_54505_58244 (
    .I(net_54505),
    .O(net_58244)
  );
  Odrv4 odrv_14_15_54507_54291 (
    .I(net_54507),
    .O(net_54291)
  );
  Odrv4 odrv_14_15_54509_54642 (
    .I(net_54509),
    .O(net_54642)
  );
  Odrv4 odrv_14_16_54626_54406 (
    .I(net_54626),
    .O(net_54406)
  );
  Odrv4 odrv_14_16_54629_54412 (
    .I(net_54629),
    .O(net_54412)
  );
  Odrv4 odrv_14_17_54753_54537 (
    .I(net_54753),
    .O(net_54537)
  );
  Odrv4 odrv_14_18_54875_58846 (
    .I(net_54875),
    .O(net_58846)
  );
  Odrv4 odrv_14_18_54875_58853 (
    .I(net_54875),
    .O(net_58853)
  );
  Odrv4 odrv_14_18_54878_55011 (
    .I(net_54878),
    .O(net_55011)
  );
  Odrv4 odrv_14_20_55122_58973 (
    .I(net_55122),
    .O(net_58973)
  );
  Odrv4 odrv_14_20_55122_59084 (
    .I(net_55122),
    .O(net_59084)
  );
  Odrv4 odrv_14_20_55124_55020 (
    .I(net_55124),
    .O(net_55020)
  );
  Odrv4 odrv_14_26_55859_59709 (
    .I(net_55859),
    .O(net_59709)
  );
  Odrv4 odrv_14_27_55979_59842 (
    .I(net_55979),
    .O(net_59842)
  );
  Odrv4 odrv_14_28_56102_52407 (
    .I(net_56102),
    .O(net_52407)
  );
  Odrv4 odrv_14_28_56102_56245 (
    .I(net_56102),
    .O(net_56245)
  );
  Odrv4 odrv_14_2_52872_56870 (
    .I(net_52872),
    .O(net_56870)
  );
  Odrv12 odrv_14_2_52873_56584 (
    .I(net_52873),
    .O(net_56584)
  );
  Odrv4 odrv_14_7_53524_53547 (
    .I(net_53524),
    .O(net_53547)
  );
  Odrv4 odrv_14_8_53645_57495 (
    .I(net_53645),
    .O(net_57495)
  );
  Odrv4 odrv_14_8_53645_57616 (
    .I(net_53645),
    .O(net_57616)
  );
  Odrv4 odrv_14_8_53646_57259 (
    .I(net_53646),
    .O(net_57259)
  );
  Odrv4 odrv_15_10_57719_57863 (
    .I(net_57719),
    .O(net_57863)
  );
  Odrv4 odrv_15_10_57721_54022 (
    .I(net_57721),
    .O(net_54022)
  );
  Odrv4 odrv_15_10_57721_57742 (
    .I(net_57721),
    .O(net_57742)
  );
  Odrv4 odrv_15_10_57721_57868 (
    .I(net_57721),
    .O(net_57868)
  );
  Odrv4 odrv_15_10_57721_61333 (
    .I(net_57721),
    .O(net_61333)
  );
  Odrv4 odrv_15_10_57721_61692 (
    .I(net_57721),
    .O(net_61692)
  );
  Odrv4 odrv_15_10_57721_61699 (
    .I(net_57721),
    .O(net_61699)
  );
  Odrv4 odrv_15_10_57722_57870 (
    .I(net_57722),
    .O(net_57870)
  );
  Odrv12 odrv_15_10_57723_60943 (
    .I(net_57723),
    .O(net_60943)
  );
  Odrv4 odrv_15_11_57843_57978 (
    .I(net_57843),
    .O(net_57978)
  );
  Odrv4 odrv_15_11_57845_61696 (
    .I(net_57845),
    .O(net_61696)
  );
  Odrv4 odrv_15_13_58086_62051 (
    .I(net_58086),
    .O(net_62051)
  );
  Odrv4 odrv_15_13_58087_58230 (
    .I(net_58087),
    .O(net_58230)
  );
  Odrv4 odrv_15_13_58087_61824 (
    .I(net_58087),
    .O(net_61824)
  );
  Odrv4 odrv_15_13_58088_62057 (
    .I(net_58088),
    .O(net_62057)
  );
  Odrv4 odrv_15_13_58091_62053 (
    .I(net_58091),
    .O(net_62053)
  );
  Odrv4 odrv_15_13_58092_58222 (
    .I(net_58092),
    .O(net_58222)
  );
  Odrv4 odrv_15_13_58092_61818 (
    .I(net_58092),
    .O(net_61818)
  );
  Odrv4 odrv_15_14_58210_61947 (
    .I(net_58210),
    .O(net_61947)
  );
  Odrv4 odrv_15_14_58210_62178 (
    .I(net_58210),
    .O(net_62178)
  );
  Odrv4 odrv_15_14_58211_57992 (
    .I(net_58211),
    .O(net_57992)
  );
  Odrv4 odrv_15_14_58212_61823 (
    .I(net_58212),
    .O(net_61823)
  );
  Odrv4 odrv_15_14_58213_62184 (
    .I(net_58213),
    .O(net_62184)
  );
  Odrv4 odrv_15_14_58215_58110 (
    .I(net_58215),
    .O(net_58110)
  );
  Odrv4 odrv_15_14_58216_58349 (
    .I(net_58216),
    .O(net_58349)
  );
  Odrv4 odrv_15_14_58216_61943 (
    .I(net_58216),
    .O(net_61943)
  );
  Odrv4 odrv_15_15_58334_62303 (
    .I(net_58334),
    .O(net_62303)
  );
  Odrv4 odrv_15_15_58335_58243 (
    .I(net_58335),
    .O(net_58243)
  );
  Odrv4 odrv_15_15_58336_62307 (
    .I(net_58336),
    .O(net_62307)
  );
  Odrv4 odrv_15_15_58338_62064 (
    .I(net_58338),
    .O(net_62064)
  );
  Odrv4 odrv_15_16_58455_58234 (
    .I(net_58455),
    .O(net_58234)
  );
  Odrv4 odrv_15_16_58458_58240 (
    .I(net_58458),
    .O(net_58240)
  );
  Odrv4 odrv_15_16_58459_62071 (
    .I(net_58459),
    .O(net_62071)
  );
  Odrv4 odrv_15_16_58460_54764 (
    .I(net_58460),
    .O(net_54764)
  );
  Odrv4 odrv_15_16_58462_58358 (
    .I(net_58462),
    .O(net_58358)
  );
  Odrv4 odrv_15_17_58579_58359 (
    .I(net_58579),
    .O(net_58359)
  );
  Odrv4 odrv_15_17_58581_58489 (
    .I(net_58581),
    .O(net_58489)
  );
  Odrv4 odrv_15_17_58583_58367 (
    .I(net_58583),
    .O(net_58367)
  );
  Odrv4 odrv_15_17_58584_54889 (
    .I(net_58584),
    .O(net_54889)
  );
  Odrv4 odrv_15_18_58701_62666 (
    .I(net_58701),
    .O(net_62666)
  );
  Odrv4 odrv_15_18_58707_58837 (
    .I(net_58707),
    .O(net_58837)
  );
  Odrv4 odrv_15_19_58827_51303 (
    .I(net_58827),
    .O(net_51303)
  );
  Odrv4 odrv_15_19_58827_58609 (
    .I(net_58827),
    .O(net_58609)
  );
  Odrv4 odrv_15_19_58827_58735 (
    .I(net_58827),
    .O(net_58735)
  );
  Odrv4 odrv_15_19_58827_58962 (
    .I(net_58827),
    .O(net_58962)
  );
  Odrv4 odrv_15_19_58827_62438 (
    .I(net_58827),
    .O(net_62438)
  );
  Odrv4 odrv_15_19_58827_62566 (
    .I(net_58827),
    .O(net_62566)
  );
  Odrv4 odrv_15_19_58827_62797 (
    .I(net_58827),
    .O(net_62797)
  );
  Odrv4 odrv_15_20_58947_58726 (
    .I(net_58947),
    .O(net_58726)
  );
  Odrv4 odrv_15_20_58947_58852 (
    .I(net_58947),
    .O(net_58852)
  );
  Odrv12 odrv_15_20_58947_61435 (
    .I(net_58947),
    .O(net_61435)
  );
  Odrv4 odrv_15_20_58947_62555 (
    .I(net_58947),
    .O(net_62555)
  );
  Odrv4 odrv_15_20_58953_51432 (
    .I(net_58953),
    .O(net_51432)
  );
  Odrv4 odrv_15_20_58954_55260 (
    .I(net_58954),
    .O(net_55260)
  );
  Odrv4 odrv_15_20_58954_58850 (
    .I(net_58954),
    .O(net_58850)
  );
  Odrv4 odrv_15_21_59076_51555 (
    .I(net_59076),
    .O(net_51555)
  );
  Odrv4 odrv_15_21_59076_55381 (
    .I(net_59076),
    .O(net_55381)
  );
  Odrv4 odrv_15_21_59076_58971 (
    .I(net_59076),
    .O(net_58971)
  );
  Odrv4 odrv_15_21_59076_59206 (
    .I(net_59076),
    .O(net_59206)
  );
  Odrv4 odrv_15_21_59076_62802 (
    .I(net_59076),
    .O(net_62802)
  );
  Odrv4 odrv_15_22_59197_58980 (
    .I(net_59197),
    .O(net_58980)
  );
  Odrv4 odrv_15_22_59197_59218 (
    .I(net_59197),
    .O(net_59218)
  );
  Odrv4 odrv_15_23_59321_51799 (
    .I(net_59321),
    .O(net_51799)
  );
  Odrv4 odrv_15_23_59321_59105 (
    .I(net_59321),
    .O(net_59105)
  );
  Odrv4 odrv_15_23_59323_59219 (
    .I(net_59323),
    .O(net_59219)
  );
  Odrv4 odrv_15_25_59567_59351 (
    .I(net_59567),
    .O(net_59351)
  );
  Odrv4 odrv_15_25_59567_59589 (
    .I(net_59567),
    .O(net_59589)
  );
  Odrv4 odrv_15_25_59567_63180 (
    .I(net_59567),
    .O(net_63180)
  );
  Odrv4 odrv_15_25_59567_63418 (
    .I(net_59567),
    .O(net_63418)
  );
  Odrv4 odrv_15_27_59813_59597 (
    .I(net_59813),
    .O(net_59597)
  );
  Odrv4 odrv_15_28_59932_59838 (
    .I(net_59932),
    .O(net_59838)
  );
  Odrv4 odrv_15_28_59938_52408 (
    .I(net_59938),
    .O(net_52408)
  );
  Odrv4 odrv_15_28_59938_56244 (
    .I(net_59938),
    .O(net_56244)
  );
  Odrv4 odrv_15_29_60061_63914 (
    .I(net_60061),
    .O(net_63914)
  );
  Odrv4 odrv_15_2_56700_56732 (
    .I(net_56700),
    .O(net_56732)
  );
  Odrv4 odrv_15_3_56861_60840 (
    .I(net_56861),
    .O(net_60840)
  );
  Odrv4 odrv_15_6_57227_49700 (
    .I(net_57227),
    .O(net_49700)
  );
  Odrv4 odrv_15_6_57227_60965 (
    .I(net_57227),
    .O(net_60965)
  );
  Odrv4 odrv_15_6_57227_61203 (
    .I(net_57227),
    .O(net_61203)
  );
  Odrv4 odrv_15_8_57471_53786 (
    .I(net_57471),
    .O(net_53786)
  );
  Odrv4 odrv_15_8_57471_61207 (
    .I(net_57471),
    .O(net_61207)
  );
  Odrv4 odrv_15_9_57601_57625 (
    .I(net_57601),
    .O(net_57625)
  );
  Odrv4 odrv_15_9_57601_57751 (
    .I(net_57601),
    .O(net_57751)
  );
  Odrv12 odrv_15_9_57601_60942 (
    .I(net_57601),
    .O(net_60942)
  );
  Odrv4 odrv_16_12_61793_61826 (
    .I(net_61793),
    .O(net_61826)
  );
  Odrv4 odrv_16_12_61793_65759 (
    .I(net_61793),
    .O(net_65759)
  );
  Odrv4 odrv_16_12_61794_65658 (
    .I(net_61794),
    .O(net_65658)
  );
  Odrv4 odrv_16_12_61794_65763 (
    .I(net_61794),
    .O(net_65763)
  );
  Odrv4 odrv_16_12_61797_54275 (
    .I(net_61797),
    .O(net_54275)
  );
  Odrv4 odrv_16_12_61798_61946 (
    .I(net_61798),
    .O(net_61946)
  );
  Odrv4 odrv_16_12_61799_61929 (
    .I(net_61799),
    .O(net_61929)
  );
  Odrv4 odrv_16_13_61918_65888 (
    .I(net_61918),
    .O(net_65888)
  );
  Odrv4 odrv_16_14_62046_61942 (
    .I(net_62046),
    .O(net_61942)
  );
  Odrv4 odrv_16_15_62164_65903 (
    .I(net_62164),
    .O(net_65903)
  );
  Odrv4 odrv_16_15_62164_66134 (
    .I(net_62164),
    .O(net_66134)
  );
  Odrv4 odrv_16_15_62166_61949 (
    .I(net_62166),
    .O(net_61949)
  );
  Odrv4 odrv_16_15_62167_62189 (
    .I(net_62167),
    .O(net_62189)
  );
  Odrv4 odrv_16_15_62167_66130 (
    .I(net_62167),
    .O(net_66130)
  );
  Odrv4 odrv_16_15_62168_62298 (
    .I(net_62168),
    .O(net_62298)
  );
  Odrv4 odrv_16_15_62169_65897 (
    .I(net_62169),
    .O(net_65897)
  );
  Odrv4 odrv_16_16_62286_62066 (
    .I(net_62286),
    .O(net_62066)
  );
  Odrv4 odrv_16_16_62286_62320 (
    .I(net_62286),
    .O(net_62320)
  );
  Odrv4 odrv_16_16_62286_66024 (
    .I(net_62286),
    .O(net_66024)
  );
  Odrv4 odrv_16_16_62286_66255 (
    .I(net_62286),
    .O(net_66255)
  );
  Odrv4 odrv_16_18_62533_66503 (
    .I(net_62533),
    .O(net_66503)
  );
  Odrv4 odrv_16_28_63765_63548 (
    .I(net_63765),
    .O(net_63548)
  );
  Odrv4 odrv_16_2_60529_60710 (
    .I(net_60529),
    .O(net_60710)
  );
  Odrv4 odrv_16_2_60530_64410 (
    .I(net_60530),
    .O(net_64410)
  );
  Odrv4 odrv_16_9_61426_61571 (
    .I(net_61426),
    .O(net_61571)
  );
  Odrv4 odrv_16_9_61430_61579 (
    .I(net_61430),
    .O(net_61579)
  );
  Odrv12 odrv_16_9_61431_64773 (
    .I(net_61431),
    .O(net_64773)
  );
  Odrv4 odrv_17_0_64354_64390 (
    .I(net_64354),
    .O(net_64390)
  );
  Odrv12 odrv_17_0_64354_68077 (
    .I(net_64354),
    .O(net_68077)
  );
  Odrv4 odrv_17_0_64355_64392 (
    .I(net_64355),
    .O(net_64392)
  );
  Odrv4 odrv_17_12_65625_65768 (
    .I(net_65625),
    .O(net_65768)
  );
  Odrv4 odrv_17_13_65753_69606 (
    .I(net_65753),
    .O(net_69606)
  );
  Odrv4 odrv_17_14_65875_69727 (
    .I(net_65875),
    .O(net_69727)
  );
  Odrv4 odrv_17_15_65996_69967 (
    .I(net_65996),
    .O(net_69967)
  );
  Odrv4 odrv_17_16_66123_62428 (
    .I(net_66123),
    .O(net_62428)
  );
  Odrv4 odrv_17_16_66123_66256 (
    .I(net_66123),
    .O(net_66256)
  );
  Odrv4 odrv_17_17_66240_70209 (
    .I(net_66240),
    .O(net_70209)
  );
  Odrv4 odrv_17_17_66244_70207 (
    .I(net_66244),
    .O(net_70207)
  );
  Odrv4 odrv_17_17_66246_66379 (
    .I(net_66246),
    .O(net_66379)
  );
  Odrv4 odrv_17_18_66365_66500 (
    .I(net_66365),
    .O(net_66500)
  );
  Odrv4 odrv_17_18_66368_58847 (
    .I(net_66368),
    .O(net_58847)
  );
  Odrv12 odrv_17_18_66368_62662 (
    .I(net_66368),
    .O(net_62662)
  );
  Odrv4 odrv_17_18_66368_66498 (
    .I(net_66368),
    .O(net_66498)
  );
  Odrv4 odrv_17_18_66368_66517 (
    .I(net_66368),
    .O(net_66517)
  );
  Odrv4 odrv_17_18_66368_70349 (
    .I(net_66368),
    .O(net_70349)
  );
  Odrv4 odrv_17_18_66369_66502 (
    .I(net_66369),
    .O(net_66502)
  );
  Odrv4 odrv_17_19_66489_62789 (
    .I(net_66489),
    .O(net_62789)
  );
  Odrv4 odrv_17_19_66489_70461 (
    .I(net_66489),
    .O(net_70461)
  );
  Odrv4 odrv_17_19_66491_70344 (
    .I(net_66491),
    .O(net_70344)
  );
  Odrv4 odrv_17_20_66609_66515 (
    .I(net_66609),
    .O(net_66515)
  );
  Odrv4 odrv_17_21_66736_70350 (
    .I(net_66736),
    .O(net_70350)
  );
  Odrv4 odrv_17_29_67720_67868 (
    .I(net_67720),
    .O(net_67868)
  );
  Odrv4 odrv_17_29_67721_71574 (
    .I(net_67721),
    .O(net_71574)
  );
  Odrv4 odrv_17_29_67722_71704 (
    .I(net_67722),
    .O(net_71704)
  );
  Odrv4 odrv_17_31_67961_67748 (
    .I(net_67961),
    .O(net_67748)
  );
  Odrv4 odrv_17_9_65256_65290 (
    .I(net_65256),
    .O(net_65290)
  );
  Odrv4 odrv_18_0_68185_68093 (
    .I(net_68185),
    .O(net_68093)
  );
  Odrv4 odrv_18_10_69212_61687 (
    .I(net_69212),
    .O(net_61687)
  );
  Odrv4 odrv_18_10_69212_69120 (
    .I(net_69212),
    .O(net_69120)
  );
  Odrv4 odrv_18_10_69212_69347 (
    .I(net_69212),
    .O(net_69347)
  );
  Odrv4 odrv_18_10_69212_73183 (
    .I(net_69212),
    .O(net_73183)
  );
  Odrv4 odrv_18_12_69458_73429 (
    .I(net_69458),
    .O(net_73429)
  );
  Odrv4 odrv_18_12_69461_69591 (
    .I(net_69461),
    .O(net_69591)
  );
  Odrv4 odrv_18_12_69462_65767 (
    .I(net_69462),
    .O(net_65767)
  );
  Odrv4 odrv_18_13_69578_73544 (
    .I(net_69578),
    .O(net_73544)
  );
  Odrv4 odrv_18_13_69580_73550 (
    .I(net_69580),
    .O(net_73550)
  );
  Odrv4 odrv_18_13_69581_69716 (
    .I(net_69581),
    .O(net_69716)
  );
  Odrv4 odrv_18_13_69582_73554 (
    .I(net_69582),
    .O(net_73554)
  );
  Odrv4 odrv_18_13_69583_65886 (
    .I(net_69583),
    .O(net_65886)
  );
  Odrv12 odrv_18_13_69584_65878 (
    .I(net_69584),
    .O(net_65878)
  );
  Odrv4 odrv_18_13_69585_69718 (
    .I(net_69585),
    .O(net_69718)
  );
  Odrv4 odrv_18_14_69701_73667 (
    .I(net_69701),
    .O(net_73667)
  );
  Odrv4 odrv_18_14_69703_69847 (
    .I(net_69703),
    .O(net_69847)
  );
  Odrv4 odrv_18_14_69704_73675 (
    .I(net_69704),
    .O(net_73675)
  );
  Odrv4 odrv_18_14_69706_73669 (
    .I(net_69706),
    .O(net_73669)
  );
  Odrv4 odrv_18_15_69824_73790 (
    .I(net_69824),
    .O(net_73790)
  );
  Odrv4 odrv_18_15_69826_69970 (
    .I(net_69826),
    .O(net_69970)
  );
  Odrv4 odrv_18_15_69827_73439 (
    .I(net_69827),
    .O(net_73439)
  );
  Odrv4 odrv_18_15_69828_62304 (
    .I(net_69828),
    .O(net_62304)
  );
  Odrv4 odrv_18_15_69829_73443 (
    .I(net_69829),
    .O(net_73443)
  );
  Odrv4 odrv_18_15_69830_62308 (
    .I(net_69830),
    .O(net_62308)
  );
  Odrv4 odrv_18_15_69831_69964 (
    .I(net_69831),
    .O(net_69964)
  );
  Odrv4 odrv_18_16_69949_70093 (
    .I(net_69949),
    .O(net_70093)
  );
  Odrv4 odrv_18_16_69949_73560 (
    .I(net_69949),
    .O(net_73560)
  );
  Odrv4 odrv_18_16_69949_73919 (
    .I(net_69949),
    .O(net_73919)
  );
  Odrv4 odrv_18_16_69949_73926 (
    .I(net_69949),
    .O(net_73926)
  );
  Odrv4 odrv_18_17_70070_74036 (
    .I(net_70070),
    .O(net_74036)
  );
  Odrv4 odrv_18_17_70071_74040 (
    .I(net_70071),
    .O(net_74040)
  );
  Odrv4 odrv_18_17_70072_74042 (
    .I(net_70072),
    .O(net_74042)
  );
  Odrv4 odrv_18_17_70073_62548 (
    .I(net_70073),
    .O(net_62548)
  );
  Odrv4 odrv_18_17_70074_74046 (
    .I(net_70074),
    .O(net_74046)
  );
  Odrv4 odrv_18_17_70075_74038 (
    .I(net_70075),
    .O(net_74038)
  );
  Odrv4 odrv_18_17_70076_70206 (
    .I(net_70076),
    .O(net_70206)
  );
  Odrv4 odrv_18_17_70077_66382 (
    .I(net_70077),
    .O(net_66382)
  );
  Odrv4 odrv_18_18_70195_74165 (
    .I(net_70195),
    .O(net_74165)
  );
  Odrv4 odrv_18_18_70199_70329 (
    .I(net_70199),
    .O(net_70329)
  );
  Odrv4 odrv_18_18_70200_66505 (
    .I(net_70200),
    .O(net_66505)
  );
  Odrv4 odrv_18_20_70446_74300 (
    .I(net_70446),
    .O(net_74300)
  );
  Odrv4 odrv_18_31_71794_71575 (
    .I(net_71794),
    .O(net_71575)
  );
  Odrv4 odrv_18_31_71794_75655 (
    .I(net_71794),
    .O(net_75655)
  );
  Odrv4 odrv_18_31_71795_71577 (
    .I(net_71795),
    .O(net_71577)
  );
  Odrv4 odrv_18_5_68599_61076 (
    .I(net_68599),
    .O(net_61076)
  );
  Odrv4 odrv_18_6_68718_72687 (
    .I(net_68718),
    .O(net_72687)
  );
  Odrv4 odrv_18_6_68722_72685 (
    .I(net_68722),
    .O(net_72685)
  );
  Odrv4 odrv_18_6_68723_61201 (
    .I(net_68723),
    .O(net_61201)
  );
  Odrv4 odrv_18_6_68724_65029 (
    .I(net_68724),
    .O(net_65029)
  );
  Odrv4 odrv_19_13_73409_77101 (
    .I(net_73409),
    .O(net_77101)
  );
  Odrv4 odrv_19_13_73413_69713 (
    .I(net_73413),
    .O(net_69713)
  );
  Odrv4 odrv_19_13_73415_65893 (
    .I(net_73415),
    .O(net_65893)
  );
  Odrv4 odrv_19_14_73532_73674 (
    .I(net_73532),
    .O(net_73674)
  );
  Odrv4 odrv_19_14_73533_76911 (
    .I(net_73533),
    .O(net_76911)
  );
  Odrv4 odrv_19_14_73535_76915 (
    .I(net_73535),
    .O(net_76915)
  );
  Odrv4 odrv_19_14_73536_77220 (
    .I(net_73536),
    .O(net_77220)
  );
  Odrv4 odrv_19_14_73539_77226 (
    .I(net_73539),
    .O(net_77226)
  );
  Odrv4 odrv_19_15_73659_66135 (
    .I(net_73659),
    .O(net_66135)
  );
  Odrv4 odrv_19_15_73661_77114 (
    .I(net_73661),
    .O(net_77114)
  );
  Odrv4 odrv_19_15_73662_73795 (
    .I(net_73662),
    .O(net_73795)
  );
  Odrv4 odrv_19_16_73779_77222 (
    .I(net_73779),
    .O(net_77222)
  );
  Odrv4 odrv_19_16_73781_73563 (
    .I(net_73781),
    .O(net_73563)
  );
  Odrv4 odrv_19_16_73783_70086 (
    .I(net_73783),
    .O(net_70086)
  );
  Odrv4 odrv_19_16_73785_73681 (
    .I(net_73785),
    .O(net_73681)
  );
  Odrv4 odrv_19_17_73901_77509 (
    .I(net_73901),
    .O(net_77509)
  );
  Odrv4 odrv_19_17_73902_77513 (
    .I(net_73902),
    .O(net_77513)
  );
  Odrv4 odrv_19_17_73903_77219 (
    .I(net_73903),
    .O(net_77219)
  );
  Odrv4 odrv_19_17_73907_70211 (
    .I(net_73907),
    .O(net_70211)
  );
  Odrv4 odrv_19_18_74028_74175 (
    .I(net_74028),
    .O(net_74175)
  );
  Odrv4 odrv_20_10_76651_80206 (
    .I(net_76651),
    .O(net_80206)
  );
  Odrv4 odrv_20_10_76654_76508 (
    .I(net_76654),
    .O(net_76508)
  );
  Odrv4 odrv_20_10_76656_80208 (
    .I(net_76656),
    .O(net_80208)
  );
  Odrv4 odrv_20_10_76658_76800 (
    .I(net_76658),
    .O(net_76800)
  );
  Odrv4 odrv_20_10_76658_76817 (
    .I(net_76658),
    .O(net_76817)
  );
  Odrv12 odrv_20_10_76658_79589 (
    .I(net_76658),
    .O(net_79589)
  );
  Odrv4 odrv_20_10_76658_79975 (
    .I(net_76658),
    .O(net_79975)
  );
  Odrv4 odrv_20_10_76658_80101 (
    .I(net_76658),
    .O(net_80101)
  );
  Odrv4 odrv_20_10_76658_80229 (
    .I(net_76658),
    .O(net_80229)
  );
  Odrv4 odrv_20_13_76958_73546 (
    .I(net_76958),
    .O(net_73546)
  );
  Odrv4 odrv_20_13_76959_69714 (
    .I(net_76959),
    .O(net_69714)
  );
  Odrv4 odrv_20_13_76960_76919 (
    .I(net_76960),
    .O(net_76919)
  );
  Odrv4 odrv_20_13_76962_69722 (
    .I(net_76962),
    .O(net_69722)
  );
  Odrv4 odrv_20_13_76963_77016 (
    .I(net_76963),
    .O(net_77016)
  );
  Odrv4 odrv_20_15_77167_77113 (
    .I(net_77167),
    .O(net_77113)
  );
  Odrv4 odrv_20_15_77168_77115 (
    .I(net_77168),
    .O(net_77115)
  );
  Odrv4 odrv_20_16_77264_77116 (
    .I(net_77264),
    .O(net_77116)
  );
  Odrv4 odrv_20_16_77264_77328 (
    .I(net_77264),
    .O(net_77328)
  );
  Odrv4 odrv_20_16_77265_77223 (
    .I(net_77265),
    .O(net_77223)
  );
  Odrv4 odrv_20_16_77265_80950 (
    .I(net_77265),
    .O(net_80950)
  );
  Odrv4 odrv_20_16_77266_77120 (
    .I(net_77266),
    .O(net_77120)
  );
  Odrv4 odrv_20_16_77266_77421 (
    .I(net_77266),
    .O(net_77421)
  );
  Odrv4 odrv_20_16_77267_77122 (
    .I(net_77267),
    .O(net_77122)
  );
  Odrv4 odrv_20_16_77267_77423 (
    .I(net_77267),
    .O(net_77423)
  );
  Odrv4 odrv_20_16_77268_77124 (
    .I(net_77268),
    .O(net_77124)
  );
  Odrv4 odrv_20_16_77268_80835 (
    .I(net_77268),
    .O(net_80835)
  );
  Odrv4 odrv_20_16_77269_77322 (
    .I(net_77269),
    .O(net_77322)
  );
  Odrv4 odrv_20_16_77270_77217 (
    .I(net_77270),
    .O(net_77217)
  );
  Odrv4 odrv_20_16_77270_80839 (
    .I(net_77270),
    .O(net_80839)
  );
  Odrv4 odrv_20_17_77365_80710 (
    .I(net_77365),
    .O(net_80710)
  );
  Odrv4 odrv_20_17_77369_80718 (
    .I(net_77369),
    .O(net_80718)
  );
  Odrv4 odrv_20_18_77472_81081 (
    .I(net_77472),
    .O(net_81081)
  );
  Odrv4 odrv_20_6_76243_79611 (
    .I(net_76243),
    .O(net_79611)
  );
  Odrv4 odrv_20_6_76245_79720 (
    .I(net_76245),
    .O(net_79720)
  );
  Odrv4 odrv_20_7_76345_76408 (
    .I(net_76345),
    .O(net_76408)
  );
  Odrv4 odrv_20_7_76345_76496 (
    .I(net_76345),
    .O(net_76496)
  );
  Odrv4 odrv_20_7_76345_79480 (
    .I(net_76345),
    .O(net_79480)
  );
  Odrv4 odrv_20_7_76345_79734 (
    .I(net_76345),
    .O(net_79734)
  );
  Odrv4 odrv_20_9_76549_79980 (
    .I(net_76549),
    .O(net_79980)
  );
  Odrv4 odrv_20_9_76550_76402 (
    .I(net_76550),
    .O(net_76402)
  );
  Odrv4 odrv_20_9_76550_79856 (
    .I(net_76550),
    .O(net_79856)
  );
  Odrv4 odrv_21_10_80072_76797 (
    .I(net_80072),
    .O(net_76797)
  );
  Odrv4 odrv_21_10_80072_79978 (
    .I(net_80072),
    .O(net_79978)
  );
  Odrv4 odrv_21_10_80072_80106 (
    .I(net_80072),
    .O(net_80106)
  );
  Odrv4 odrv_21_10_80072_80215 (
    .I(net_80072),
    .O(net_80215)
  );
  Odrv12 odrv_21_10_80072_83666 (
    .I(net_80072),
    .O(net_83666)
  );
  Odrv4 odrv_21_10_80072_84041 (
    .I(net_80072),
    .O(net_84041)
  );
  Odrv4 odrv_21_10_80075_76795 (
    .I(net_80075),
    .O(net_76795)
  );
  Odrv4 odrv_21_10_80075_80096 (
    .I(net_80075),
    .O(net_80096)
  );
  Odrv4 odrv_21_10_80075_80222 (
    .I(net_80075),
    .O(net_80222)
  );
  Odrv4 odrv_21_10_80075_83926 (
    .I(net_80075),
    .O(net_83926)
  );
  Odrv4 odrv_21_10_80075_84047 (
    .I(net_80075),
    .O(net_84047)
  );
  Odrv4 odrv_21_10_80076_84039 (
    .I(net_80076),
    .O(net_84039)
  );
  Odrv4 odrv_21_12_80322_80470 (
    .I(net_80322),
    .O(net_80470)
  );
  Odrv4 odrv_21_13_80440_80473 (
    .I(net_80440),
    .O(net_80473)
  );
  Odrv4 odrv_21_13_80443_80589 (
    .I(net_80443),
    .O(net_80589)
  );
  Odrv4 odrv_21_13_80444_84423 (
    .I(net_80444),
    .O(net_84423)
  );
  Odrv4 odrv_21_14_80563_80596 (
    .I(net_80563),
    .O(net_80596)
  );
  Odrv4 odrv_21_14_80569_80464 (
    .I(net_80569),
    .O(net_80464)
  );
  Odrv4 odrv_21_16_80813_77407 (
    .I(net_80813),
    .O(net_77407)
  );
  Odrv4 odrv_21_17_80938_74047 (
    .I(net_80938),
    .O(net_74047)
  );
  Odrv4 odrv_21_17_80938_80833 (
    .I(net_80938),
    .O(net_80833)
  );
  Odrv4 odrv_21_17_80938_81068 (
    .I(net_80938),
    .O(net_81068)
  );
  Odrv4 odrv_21_17_80938_84665 (
    .I(net_80938),
    .O(net_84665)
  );
  Odrv12 odrv_21_18_81055_70324 (
    .I(net_81055),
    .O(net_70324)
  );
  Odrv4 odrv_21_18_81057_80838 (
    .I(net_81057),
    .O(net_80838)
  );
  Odrv4 odrv_21_18_81060_80844 (
    .I(net_81060),
    .O(net_80844)
  );
  Odrv4 odrv_21_18_81062_80958 (
    .I(net_81062),
    .O(net_80958)
  );
  Odrv4 odrv_21_19_81181_80963 (
    .I(net_81181),
    .O(net_80963)
  );
  Odrv4 odrv_21_6_79582_83194 (
    .I(net_79582),
    .O(net_83194)
  );
  Odrv4 odrv_21_6_79584_72692 (
    .I(net_79584),
    .O(net_72692)
  );
  Odrv4 odrv_21_6_79584_76391 (
    .I(net_79584),
    .O(net_76391)
  );
  Odrv4 odrv_21_6_79584_79368 (
    .I(net_79584),
    .O(net_79368)
  );
  Odrv4 odrv_21_6_79584_79732 (
    .I(net_79584),
    .O(net_79732)
  );
  Odrv12 odrv_21_6_79584_82776 (
    .I(net_79584),
    .O(net_82776)
  );
  Odrv4 odrv_21_6_79584_83198 (
    .I(net_79584),
    .O(net_83198)
  );
  Odrv4 odrv_21_6_79584_83547 (
    .I(net_79584),
    .O(net_83547)
  );
  Odrv4 odrv_21_6_79584_83564 (
    .I(net_79584),
    .O(net_83564)
  );
  Odrv4 odrv_21_9_79948_83914 (
    .I(net_79948),
    .O(net_83914)
  );
  Odrv4 odrv_21_9_79950_80094 (
    .I(net_79950),
    .O(net_80094)
  );
  Odrv4 odrv_21_9_79950_80095 (
    .I(net_79950),
    .O(net_80095)
  );
  Odrv12 odrv_21_9_79950_83667 (
    .I(net_79950),
    .O(net_83667)
  );
  Odrv4 odrv_21_9_79954_76699 (
    .I(net_79954),
    .O(net_76699)
  );
  Odrv4 odrv_22_13_84276_77110 (
    .I(net_84276),
    .O(net_77110)
  );
  Odrv4 odrv_22_14_84397_77208 (
    .I(net_84397),
    .O(net_77208)
  );
  Odrv4 odrv_22_15_84519_84664 (
    .I(net_84519),
    .O(net_84664)
  );
  Odrv4 odrv_22_15_84519_88496 (
    .I(net_84519),
    .O(net_88496)
  );
  Odrv4 odrv_22_17_84764_84544 (
    .I(net_84764),
    .O(net_84544)
  );
  Odrv4 odrv_22_17_84764_84798 (
    .I(net_84764),
    .O(net_84798)
  );
  Odrv4 odrv_22_17_84764_84907 (
    .I(net_84764),
    .O(net_84907)
  );
  Odrv4 odrv_22_17_84764_88374 (
    .I(net_84764),
    .O(net_88374)
  );
  Odrv4 odrv_22_17_84765_77510 (
    .I(net_84765),
    .O(net_77510)
  );
  Odrv4 odrv_22_17_84765_88376 (
    .I(net_84765),
    .O(net_88376)
  );
  Odrv4 odrv_22_17_84766_77514 (
    .I(net_84766),
    .O(net_77514)
  );
  Odrv4 odrv_22_17_84766_84548 (
    .I(net_84766),
    .O(net_84548)
  );
  Odrv4 odrv_22_17_84766_84901 (
    .I(net_84766),
    .O(net_84901)
  );
  Odrv4 odrv_22_17_84767_77516 (
    .I(net_84767),
    .O(net_77516)
  );
  Odrv4 odrv_22_17_84767_84550 (
    .I(net_84767),
    .O(net_84550)
  );
  Odrv4 odrv_22_17_84767_88739 (
    .I(net_84767),
    .O(net_88739)
  );
  Odrv4 odrv_22_17_84768_77518 (
    .I(net_84768),
    .O(net_77518)
  );
  Odrv4 odrv_22_17_84768_88382 (
    .I(net_84768),
    .O(net_88382)
  );
  Odrv4 odrv_22_17_84769_84792 (
    .I(net_84769),
    .O(net_84792)
  );
  Odrv4 odrv_22_17_84769_84899 (
    .I(net_84769),
    .O(net_84899)
  );
  Odrv4 odrv_22_17_84770_77512 (
    .I(net_84770),
    .O(net_77512)
  );
  Odrv4 odrv_22_17_84770_84666 (
    .I(net_84770),
    .O(net_84666)
  );
  Odrv4 odrv_22_17_84770_84903 (
    .I(net_84770),
    .O(net_84903)
  );
  Odrv4 odrv_23_9_87617_87513 (
    .I(net_87617),
    .O(net_87513)
  );
  Odrv4 odrv_2_19_9360_13619 (
    .I(net_9360),
    .O(net_13619)
  );
  Odrv4 odrv_2_8_7750_12035 (
    .I(net_7750),
    .O(net_12035)
  );
  Odrv4 odrv_2_8_7750_1816 (
    .I(net_7750),
    .O(net_1816)
  );
  Odrv4 odrv_3_13_12753_12886 (
    .I(net_12753),
    .O(net_12886)
  );
  Odrv12 odrv_3_13_12753_16095 (
    .I(net_12753),
    .O(net_16095)
  );
  Odrv4 odrv_3_13_12753_2864 (
    .I(net_12753),
    .O(net_2864)
  );
  Odrv4 odrv_3_7_12015_12039 (
    .I(net_12015),
    .O(net_12039)
  );
  Odrv4 odrv_4_12_16456_20426 (
    .I(net_16456),
    .O(net_20426)
  );
  Odrv4 odrv_4_13_16582_16366 (
    .I(net_16582),
    .O(net_16366)
  );
  Odrv4 odrv_4_18_17194_20805 (
    .I(net_17194),
    .O(net_20805)
  );
  Odrv4 odrv_4_18_17194_20933 (
    .I(net_17194),
    .O(net_20933)
  );
  Odrv4 odrv_4_18_17194_21164 (
    .I(net_17194),
    .O(net_21164)
  );
  Odrv4 odrv_4_18_17194_21171 (
    .I(net_17194),
    .O(net_21171)
  );
  Odrv4 odrv_4_18_17199_17095 (
    .I(net_17199),
    .O(net_17095)
  );
  Odrv4 odrv_5_12_20287_24257 (
    .I(net_20287),
    .O(net_24257)
  );
  Odrv4 odrv_5_20_21271_25241 (
    .I(net_21271),
    .O(net_25241)
  );
  Odrv4 odrv_5_5_19424_23161 (
    .I(net_19424),
    .O(net_23161)
  );
  Odrv4 odrv_5_5_19424_23390 (
    .I(net_19424),
    .O(net_23390)
  );
  Odrv4 odrv_6_0_22846_22900 (
    .I(net_22846),
    .O(net_22900)
  );
  Odrv12 odrv_6_0_22847_26571 (
    .I(net_22847),
    .O(net_26571)
  );
  Odrv4 odrv_7_0_26625_26691 (
    .I(net_26625),
    .O(net_26691)
  );
  Odrv4 odrv_7_12_27690_31284 (
    .I(net_27690),
    .O(net_31284)
  );
  Odrv4 odrv_8_10_30908_24008 (
    .I(net_30908),
    .O(net_24008)
  );
  Odrv4 odrv_8_10_30908_27633 (
    .I(net_30908),
    .O(net_27633)
  );
  Odrv4 odrv_8_10_30908_31041 (
    .I(net_30908),
    .O(net_31041)
  );
  Odrv12 odrv_8_10_30908_34250 (
    .I(net_30908),
    .O(net_34250)
  );
  Odrv4 odrv_8_12_31148_30928 (
    .I(net_31148),
    .O(net_30928)
  );
  Odrv4 odrv_8_12_31148_35117 (
    .I(net_31148),
    .O(net_35117)
  );
  Odrv4 odrv_8_17_31767_28343 (
    .I(net_31767),
    .O(net_28343)
  );
  Odrv4 odrv_8_17_31767_35747 (
    .I(net_31767),
    .O(net_35747)
  );
  Odrv4 odrv_8_23_32505_32527 (
    .I(net_32505),
    .O(net_32527)
  );
  Odrv4 odrv_8_25_32752_32775 (
    .I(net_32752),
    .O(net_32775)
  );
  Odrv4 odrv_8_25_32752_32882 (
    .I(net_32752),
    .O(net_32882)
  );
  Odrv4 odrv_8_25_32752_32901 (
    .I(net_32752),
    .O(net_32901)
  );
  Odrv4 odrv_8_25_32752_36605 (
    .I(net_32752),
    .O(net_36605)
  );
  Odrv4 odrv_8_2_29885_29936 (
    .I(net_29885),
    .O(net_29936)
  );
  Odrv4 odrv_8_2_29886_26813 (
    .I(net_29886),
    .O(net_26813)
  );
  Odrv4 odrv_8_2_29888_30057 (
    .I(net_29888),
    .O(net_30057)
  );
  Odrv4 odrv_8_31_33486_33556 (
    .I(net_33486),
    .O(net_33556)
  );
  Odrv4 odrv_8_31_33486_37347 (
    .I(net_33486),
    .O(net_37347)
  );
  Odrv4 odrv_8_3_30041_30184 (
    .I(net_30041),
    .O(net_30184)
  );
  Odrv4 odrv_8_3_30041_33774 (
    .I(net_30041),
    .O(net_33774)
  );
  Odrv4 odrv_8_3_30047_26919 (
    .I(net_30047),
    .O(net_26919)
  );
  Odrv4 odrv_8_4_30164_27015 (
    .I(net_30164),
    .O(net_27015)
  );
  Odrv4 odrv_8_4_30164_30198 (
    .I(net_30164),
    .O(net_30198)
  );
  Odrv4 odrv_8_4_30164_30307 (
    .I(net_30164),
    .O(net_30307)
  );
  Odrv12 odrv_8_4_30164_33722 (
    .I(net_30164),
    .O(net_33722)
  );
  Odrv4 odrv_8_4_30164_33768 (
    .I(net_30164),
    .O(net_33768)
  );
  Odrv4 odrv_8_4_30164_34028 (
    .I(net_30164),
    .O(net_34028)
  );
  Odrv4 odrv_8_4_30164_34133 (
    .I(net_30164),
    .O(net_34133)
  );
  Odrv4 odrv_9_10_34733_38702 (
    .I(net_34733),
    .O(net_38702)
  );
  Odrv4 odrv_9_10_34736_38715 (
    .I(net_34736),
    .O(net_38715)
  );
  Odrv4 odrv_9_10_34738_34868 (
    .I(net_34738),
    .O(net_34868)
  );
  Odrv4 odrv_9_11_34860_38823 (
    .I(net_34860),
    .O(net_38823)
  );
  Odrv4 odrv_9_12_34979_34759 (
    .I(net_34979),
    .O(net_34759)
  );
  Odrv4 odrv_9_12_34979_38589 (
    .I(net_34979),
    .O(net_38589)
  );
  Odrv4 odrv_9_12_34979_38843 (
    .I(net_34979),
    .O(net_38843)
  );
  Odrv4 odrv_9_18_35717_39686 (
    .I(net_35717),
    .O(net_39686)
  );
  Odrv4 odrv_9_18_35721_39335 (
    .I(net_35721),
    .O(net_39335)
  );
  Odrv4 odrv_9_28_36947_33252 (
    .I(net_36947),
    .O(net_33252)
  );
  Odrv4 odrv_9_28_36952_37101 (
    .I(net_36952),
    .O(net_37101)
  );
  Odrv4 odrv_9_29_37072_29568 (
    .I(net_37072),
    .O(net_29568)
  );
  Odrv4 odrv_9_4_33994_33899 (
    .I(net_33994),
    .O(net_33899)
  );
  Odrv4 odrv_9_5_34120_37860 (
    .I(net_34120),
    .O(net_37860)
  );
  Odrv4 odrv_9_8_34488_38227 (
    .I(net_34488),
    .O(net_38227)
  );
  Odrv4 odrv_9_8_34489_38229 (
    .I(net_34489),
    .O(net_38229)
  );
  Odrv4 odrv_9_8_34490_30790 (
    .I(net_34490),
    .O(net_30790)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b000001)
  ) pre_io_12_31_1 (
    .CLOCKENABLE(),
    .DIN0(net_48810),
    .DIN1(),
    .DOUT0(),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_12_31_1_dout),
    .PADOEN(io_pad_12_31_1_oe),
    .PADOUT(io_pad_12_31_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b110100)
  ) pre_io_13_31_0 (
    .CLOCKENABLE(net_56521),
    .DIN0(net_52639),
    .DIN1(net_52640),
    .DOUT0(net_56515),
    .DOUT1(),
    .INPUTCLK(net_56522),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(net_56523),
    .OUTPUTENABLE(),
    .PADIN(io_pad_13_31_0_dout),
    .PADOEN(io_pad_13_31_0_oe),
    .PADOUT(io_pad_13_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b110100)
  ) pre_io_17_0_0 (
    .CLOCKENABLE(net_68042),
    .DIN0(net_64354),
    .DIN1(net_64355),
    .DOUT0(net_68036),
    .DOUT1(),
    .INPUTCLK(net_68043),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(net_68044),
    .OUTPUTENABLE(),
    .PADIN(io_pad_17_0_0_dout),
    .PADOEN(io_pad_17_0_0_oe),
    .PADOUT(io_pad_17_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b110100)
  ) pre_io_17_31_0 (
    .CLOCKENABLE(net_71843),
    .DIN0(net_67961),
    .DIN1(),
    .DOUT0(net_71837),
    .DOUT1(),
    .INPUTCLK(net_71844),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(net_71845),
    .OUTPUTENABLE(),
    .PADIN(io_pad_17_31_0_dout),
    .PADOEN(io_pad_17_31_0_oe),
    .PADOUT(io_pad_17_31_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b110100)
  ) pre_io_18_0_0 (
    .CLOCKENABLE(net_71873),
    .DIN0(net_68185),
    .DIN1(),
    .DOUT0(net_71867),
    .DOUT1(),
    .INPUTCLK(net_71874),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(net_71875),
    .OUTPUTENABLE(),
    .PADIN(io_pad_18_0_0_dout),
    .PADOEN(io_pad_18_0_0_oe),
    .PADOUT(io_pad_18_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b110100)
  ) pre_io_18_31_1 (
    .CLOCKENABLE(net_75674),
    .DIN0(net_71794),
    .DIN1(net_71795),
    .DOUT0(net_75671),
    .DOUT1(),
    .INPUTCLK(net_75675),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(net_75676),
    .OUTPUTENABLE(),
    .PADIN(io_pad_18_31_1_dout),
    .PADOEN(io_pad_18_31_1_oe),
    .PADOUT(io_pad_18_31_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b011001)
  ) pre_io_22_0_1 (
    .CLOCKENABLE(),
    .DIN0(),
    .DIN1(),
    .DOUT0(net_86563),
    .DOUT1(),
    .INPUTCLK(),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(),
    .OUTPUTENABLE(),
    .PADIN(io_pad_22_0_1_dout),
    .PADOEN(io_pad_22_0_1_oe),
    .PADOUT(io_pad_22_0_1_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b110100)
  ) pre_io_6_0_0 (
    .CLOCKENABLE(net_26534),
    .DIN0(net_22846),
    .DIN1(net_22847),
    .DOUT0(net_26528),
    .DOUT1(),
    .INPUTCLK(net_26535),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(net_26536),
    .OUTPUTENABLE(),
    .PADIN(io_pad_6_0_0_dout),
    .PADOEN(io_pad_6_0_0_oe),
    .PADOUT(io_pad_6_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b110100)
  ) pre_io_7_0_0 (
    .CLOCKENABLE(net_29734),
    .DIN0(net_26625),
    .DIN1(),
    .DOUT0(net_29728),
    .DOUT1(),
    .INPUTCLK(net_29735),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(net_29736),
    .OUTPUTENABLE(),
    .PADIN(io_pad_7_0_0_dout),
    .PADOEN(io_pad_7_0_0_oe),
    .PADOUT(io_pad_7_0_0_din)
  );
  PRE_IO #(
    .NEG_TRIGGER(1'b0),
    .PIN_TYPE(6'b110100)
  ) pre_io_8_31_1 (
    .CLOCKENABLE(net_37366),
    .DIN0(net_33486),
    .DIN1(),
    .DOUT0(net_37363),
    .DOUT1(),
    .INPUTCLK(net_37367),
    .LATCHINPUTVALUE(),
    .OUTPUTCLK(net_37368),
    .OUTPUTENABLE(),
    .PADIN(io_pad_8_31_1_dout),
    .PADOEN(io_pad_8_31_1_oe),
    .PADOUT(io_pad_8_31_1_din)
  );
  SB_RAM40_4K ram_19_13 (
    .RCLK(net_77086),
    .RCLKE(net_77087),
    .RE(net_77088),
    .WCLK(net_77188),
    .WCLKE(net_77189),
    .WE(net_77198),
    .MASK({dangling_wire_6, dangling_wire_5, dangling_wire_4, dangling_wire_3, dangling_wire_2, dangling_wire_1, dangling_wire_15, dangling_wire_14, dangling_wire_13, dangling_wire_12, dangling_wire_11, dangling_wire_10, dangling_wire_9, dangling_wire_8, dangling_wire_7, dangling_wire_0}),
    .RADDR({dangling_wire_16, dangling_wire_18, dangling_wire_17, net_77083_cascademuxed, net_77082_cascademuxed, net_77081_cascademuxed, net_77080_cascademuxed, net_77079_cascademuxed, net_77078_cascademuxed, net_77076_cascademuxed, net_77075_cascademuxed}),
    .RDATA({net_73409, net_73410, net_73411, net_73412, net_73413, net_73414, net_73415, net_73416, net_73532, net_73533, net_73534, net_73535, net_73536, net_73537, net_73538, net_73539}),
    .WADDR({dangling_wire_19, dangling_wire_21, dangling_wire_20, net_77185_cascademuxed, net_77184_cascademuxed, net_77183_cascademuxed, net_77182_cascademuxed, net_77181_cascademuxed, net_77180_cascademuxed, net_77178_cascademuxed, net_77177_cascademuxed}),
    .WDATA({net_77094, net_77093, net_77092, net_77091, net_77090, net_77089, net_77096, net_77095, net_77197, net_77196, net_77195, net_77194, net_77193, net_77192, net_77191, net_77190})
  );
  SB_RAM40_4K ram_19_15 (
    .RCLK(net_77290),
    .RCLKE(net_77291),
    .RE(net_77292),
    .WCLK(net_77392),
    .WCLKE(net_77393),
    .WE(net_77402),
    .MASK({dangling_wire_28, dangling_wire_27, dangling_wire_26, dangling_wire_25, dangling_wire_24, dangling_wire_23, dangling_wire_37, dangling_wire_36, dangling_wire_35, dangling_wire_34, dangling_wire_33, dangling_wire_32, dangling_wire_31, dangling_wire_30, dangling_wire_29, dangling_wire_22}),
    .RADDR({dangling_wire_38, dangling_wire_40, dangling_wire_39, net_77287_cascademuxed, net_77286_cascademuxed, net_77285_cascademuxed, net_77284_cascademuxed, net_77283_cascademuxed, net_77282_cascademuxed, net_77280_cascademuxed, net_77279_cascademuxed}),
    .RDATA({net_73655, net_73656, net_73657, net_73658, net_73659, net_73660, net_73661, net_73662, net_73778, net_73779, net_73780, net_73781, net_73782, net_73783, net_73784, net_73785}),
    .WADDR({dangling_wire_41, dangling_wire_43, dangling_wire_42, net_77389_cascademuxed, net_77388_cascademuxed, net_77387_cascademuxed, net_77386_cascademuxed, net_77385_cascademuxed, net_77384_cascademuxed, net_77382_cascademuxed, net_77381_cascademuxed}),
    .WDATA({net_77298, net_77297, net_77296, net_77295, net_77294, net_77293, net_77300, net_77299, net_77401, net_77400, net_77399, net_77398, net_77397, net_77396, net_77395, net_77394})
  );
  SB_RAM40_4K ram_19_17 (
    .RCLK(net_77494),
    .RCLKE(net_77495),
    .RE(net_77496),
    .WCLK(net_77596),
    .WCLKE(net_77597),
    .WE(net_77606),
    .MASK({dangling_wire_50, dangling_wire_49, dangling_wire_48, dangling_wire_47, dangling_wire_46, dangling_wire_45, dangling_wire_59, dangling_wire_58, dangling_wire_57, dangling_wire_56, dangling_wire_55, dangling_wire_54, dangling_wire_53, dangling_wire_52, dangling_wire_51, dangling_wire_44}),
    .RADDR({dangling_wire_60, dangling_wire_62, dangling_wire_61, net_77491_cascademuxed, net_77490_cascademuxed, net_77489_cascademuxed, net_77488_cascademuxed, net_77487_cascademuxed, net_77486_cascademuxed, net_77484_cascademuxed, net_77483_cascademuxed}),
    .RDATA({net_73901, net_73902, net_73903, net_73904, net_73905, net_73906, net_73907, net_73908, net_74024, net_74025, net_74026, net_74027, net_74028, net_74029, net_74030, net_74031}),
    .WADDR({dangling_wire_63, dangling_wire_65, dangling_wire_64, net_77593_cascademuxed, net_77592_cascademuxed, net_77591_cascademuxed, net_77590_cascademuxed, net_77589_cascademuxed, net_77588_cascademuxed, net_77586_cascademuxed, net_77585_cascademuxed}),
    .WDATA({dangling_wire_66, net_77501, net_77500, net_77499, net_77498, net_77497, net_77504, net_77503, net_77605, net_77604, net_77603, net_77602, net_77601, net_77600, net_77599, net_77598})
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t1 (
    .carryinitin(),
    .carryinitout(t0)
  );
  CascadeMux t100 (
    .I(net_38393),
    .O(net_38393_cascademuxed)
  );
  LocalMux t1000 (
    .I(seg_11_23_sp4_r_v_b_19_47732),
    .O(seg_11_23_local_g3_3_47892)
  );
  Span4Mux_v4 t1001 (
    .I(seg_12_20_sp4_v_b_10_47244),
    .O(seg_11_23_sp4_r_v_b_19_47732)
  );
  Span4Mux_v4 t1002 (
    .I(seg_12_16_sp4_v_b_10_46752),
    .O(seg_12_20_sp4_v_b_10_47244)
  );
  Span4Mux_v4 t1003 (
    .I(seg_12_12_sp4_v_b_10_46260),
    .O(seg_12_16_sp4_v_b_10_46752)
  );
  Span4Mux_v4 t1004 (
    .I(seg_12_8_sp4_v_b_2_45760),
    .O(seg_12_12_sp4_v_b_10_46260)
  );
  Span4Mux_v4 t1005 (
    .I(seg_12_4_sp4_h_l_39_34133),
    .O(seg_12_8_sp4_v_b_2_45760)
  );
  LocalMux t1006 (
    .I(seg_12_28_sp4_v_b_9_48225),
    .O(seg_12_28_local_g1_1_52320)
  );
  Span4Mux_v4 t1007 (
    .I(seg_12_24_sp4_v_b_6_47732),
    .O(seg_12_28_sp4_v_b_9_48225)
  );
  Span4Mux_v4 t1008 (
    .I(seg_12_20_sp4_v_b_10_47244),
    .O(seg_12_24_sp4_v_b_6_47732)
  );
  LocalMux t1009 (
    .I(seg_14_4_sp4_h_r_29_49460),
    .O(seg_14_4_local_g2_5_57041)
  );
  CascadeMux t101 (
    .I(net_38405),
    .O(net_38405_cascademuxed)
  );
  Span4Mux_h4 t1010 (
    .I(seg_12_4_sp4_h_l_39_34133),
    .O(seg_14_4_sp4_h_r_29_49460)
  );
  LocalMux t1011 (
    .I(seg_15_16_sp4_r_v_b_5_62067),
    .O(seg_15_16_local_g1_5_62339)
  );
  Span4Mux_v4 t1012 (
    .I(seg_16_12_sp4_v_b_5_61575),
    .O(seg_15_16_sp4_r_v_b_5_62067)
  );
  Span4Mux_v4 t1013 (
    .I(seg_16_8_sp4_v_b_5_61083),
    .O(seg_16_12_sp4_v_b_5_61575)
  );
  Span4Mux_v4 t1014 (
    .I(seg_16_4_sp4_h_l_40_49460),
    .O(seg_16_8_sp4_v_b_5_61083)
  );
  Span4Mux_h4 t1015 (
    .I(seg_12_4_sp4_h_l_39_34133),
    .O(seg_16_4_sp4_h_l_40_49460)
  );
  LocalMux t1016 (
    .I(seg_19_16_sp4_h_r_42_66260),
    .O(seg_19_16_local_g2_2_77351)
  );
  Span4Mux_h4 t1017 (
    .I(seg_16_16_sp4_h_l_41_50935),
    .O(seg_19_16_sp4_h_r_42_66260)
  );
  Span4Mux_h4 t1018 (
    .I(seg_12_16_sp4_v_b_10_46752),
    .O(seg_16_16_sp4_h_l_41_50935)
  );
  LocalMux t1019 (
    .I(seg_19_16_sp4_h_r_36_66252),
    .O(seg_19_16_local_g2_4_77353)
  );
  CascadeMux t102 (
    .I(net_38411),
    .O(net_38411_cascademuxed)
  );
  Span4Mux_h4 t1020 (
    .I(seg_16_16_sp4_h_l_47_50931),
    .O(seg_19_16_sp4_h_r_36_66252)
  );
  Span4Mux_h4 t1021 (
    .I(seg_12_16_sp4_v_b_10_46752),
    .O(seg_16_16_sp4_h_l_47_50931)
  );
  LocalMux t1022 (
    .I(seg_19_18_sp4_r_v_b_26_77524),
    .O(seg_19_18_local_g0_2_77539)
  );
  Span4Mux_v4 t1023 (
    .I(seg_20_16_sp4_v_b_11_77123),
    .O(seg_19_18_sp4_r_v_b_26_77524)
  );
  Span4Mux_v4 t1024 (
    .I(seg_20_12_sp4_v_b_8_76714),
    .O(seg_20_16_sp4_v_b_11_77123)
  );
  Span4Mux_v4 t1025 (
    .I(seg_20_8_sp4_v_b_5_76301),
    .O(seg_20_12_sp4_v_b_8_76714)
  );
  Span4Mux_v4 t1026 (
    .I(seg_20_4_sp4_h_l_40_64782),
    .O(seg_20_8_sp4_v_b_5_76301)
  );
  Span4Mux_h4 t1027 (
    .I(seg_16_4_sp4_h_l_40_49460),
    .O(seg_20_4_sp4_h_l_40_64782)
  );
  LocalMux t1028 (
    .I(seg_19_18_sp4_r_v_b_29_77525),
    .O(seg_19_18_local_g1_5_77550)
  );
  Span4Mux_v4 t1029 (
    .I(seg_20_16_sp4_v_b_9_77121),
    .O(seg_19_18_sp4_r_v_b_29_77525)
  );
  CascadeMux t103 (
    .I(net_38417),
    .O(net_38417_cascademuxed)
  );
  Span4Mux_v4 t1030 (
    .I(seg_20_12_sp4_v_b_1_76705),
    .O(seg_20_16_sp4_v_b_9_77121)
  );
  Span4Mux_v4 t1031 (
    .I(seg_20_8_sp4_v_b_5_76301),
    .O(seg_20_12_sp4_v_b_1_76705)
  );
  LocalMux t1032 (
    .I(seg_6_0_span4_vert_42_22911),
    .O(seg_6_0_local_g1_2_26547)
  );
  Span4Mux_v4 t1033 (
    .I(seg_6_4_sp4_h_l_36_11775),
    .O(seg_6_0_span4_vert_42_22911)
  );
  Span4Mux_h4 t1034 (
    .I(seg_6_4_sp4_h_r_10_27015),
    .O(seg_6_4_sp4_h_l_36_11775)
  );
  LocalMux t1035 (
    .I(seg_9_27_sp4_r_v_b_16_40559),
    .O(seg_9_27_local_g3_0_40719)
  );
  Span4Mux_v4 t1036 (
    .I(seg_10_24_sp4_v_b_9_40071),
    .O(seg_9_27_sp4_r_v_b_16_40559)
  );
  Span4Mux_v4 t1037 (
    .I(seg_10_20_sp4_v_b_1_39571),
    .O(seg_10_24_sp4_v_b_9_40071)
  );
  Span4Mux_v4 t1038 (
    .I(seg_10_16_sp4_v_b_1_39079),
    .O(seg_10_20_sp4_v_b_1_39571)
  );
  Span4Mux_v4 t1039 (
    .I(seg_10_12_sp4_v_b_1_38587),
    .O(seg_10_16_sp4_v_b_1_39079)
  );
  CascadeMux t104 (
    .I(net_38423),
    .O(net_38423_cascademuxed)
  );
  Span4Mux_v4 t1040 (
    .I(seg_10_8_sp4_v_b_10_38106),
    .O(seg_10_12_sp4_v_b_1_38587)
  );
  Span4Mux_v4 t1041 (
    .I(seg_10_4_sp4_h_l_47_27015),
    .O(seg_10_8_sp4_v_b_10_38106)
  );
  LocalMux t1042 (
    .I(seg_14_9_sp4_v_b_41_53916),
    .O(seg_14_9_local_g2_1_57652)
  );
  Span4Mux_v4 t1043 (
    .I(seg_14_8_sp4_v_b_1_53419),
    .O(seg_14_9_sp4_v_b_41_53916)
  );
  Span4Mux_v4 t1044 (
    .I(seg_14_4_sp4_h_l_36_41792),
    .O(seg_14_8_sp4_v_b_1_53419)
  );
  Span4Mux_h4 t1045 (
    .I(seg_10_4_sp4_h_l_47_27015),
    .O(seg_14_4_sp4_h_l_36_41792)
  );
  LocalMux t1046 (
    .I(seg_14_9_sp4_v_b_41_53916),
    .O(seg_14_9_local_g3_1_57660)
  );
  LocalMux t1047 (
    .I(seg_14_27_sp4_v_b_18_55885),
    .O(seg_14_27_local_g0_2_59851)
  );
  Span4Mux_v4 t1048 (
    .I(seg_14_24_sp4_v_b_11_55397),
    .O(seg_14_27_sp4_v_b_18_55885)
  );
  Span4Mux_v4 t1049 (
    .I(seg_14_20_sp4_v_b_3_54897),
    .O(seg_14_24_sp4_v_b_11_55397)
  );
  CascadeMux t105 (
    .I(net_38429),
    .O(net_38429_cascademuxed)
  );
  Span4Mux_v4 t1050 (
    .I(seg_14_16_sp4_v_b_0_54404),
    .O(seg_14_20_sp4_v_b_3_54897)
  );
  Span4Mux_v4 t1051 (
    .I(seg_14_12_sp4_v_b_4_53916),
    .O(seg_14_16_sp4_v_b_0_54404)
  );
  Span4Mux_v4 t1052 (
    .I(seg_14_8_sp4_v_b_1_53419),
    .O(seg_14_12_sp4_v_b_4_53916)
  );
  LocalMux t1053 (
    .I(seg_18_0_span4_vert_42_68250),
    .O(seg_18_0_local_g0_2_71878)
  );
  Span4Mux_v4 t1054 (
    .I(seg_18_4_sp4_h_l_36_57115),
    .O(seg_18_0_span4_vert_42_68250)
  );
  Span4Mux_h4 t1055 (
    .I(seg_14_4_sp4_h_l_36_41792),
    .O(seg_18_4_sp4_h_l_36_57115)
  );
  LocalMux t1056 (
    .I(seg_18_5_sp4_v_b_43_68748),
    .O(seg_18_5_local_g2_3_72485)
  );
  Span4Mux_v4 t1057 (
    .I(seg_18_4_sp4_h_l_36_57115),
    .O(seg_18_5_sp4_v_b_43_68748)
  );
  LocalMux t1058 (
    .I(seg_9_2_sp4_v_b_27_33768),
    .O(seg_9_2_local_g2_3_37639)
  );
  LocalMux t1059 (
    .I(seg_9_12_sp4_v_b_6_34763),
    .O(seg_9_12_local_g1_6_38864)
  );
  CascadeMux t106 (
    .I(net_38645),
    .O(net_38645_cascademuxed)
  );
  Span4Mux_v4 t1060 (
    .I(seg_9_8_sp4_v_b_6_34271),
    .O(seg_9_12_sp4_v_b_6_34763)
  );
  Span4Mux_v4 t1061 (
    .I(seg_9_4_sp4_v_b_3_33768),
    .O(seg_9_8_sp4_v_b_6_34271)
  );
  LocalMux t1062 (
    .I(seg_13_31_span4_vert_18_52546),
    .O(seg_13_31_local_g1_2_56534)
  );
  Span4Mux_v4 t1063 (
    .I(seg_13_28_sp4_v_b_4_52053),
    .O(seg_13_31_span4_vert_18_52546)
  );
  Span4Mux_v4 t1064 (
    .I(seg_13_24_sp4_v_b_8_51565),
    .O(seg_13_28_sp4_v_b_4_52053)
  );
  Span4Mux_v4 t1065 (
    .I(seg_13_20_sp4_v_b_0_51065),
    .O(seg_13_24_sp4_v_b_8_51565)
  );
  Span4Mux_v4 t1066 (
    .I(seg_13_16_sp4_v_b_0_50573),
    .O(seg_13_20_sp4_v_b_0_51065)
  );
  Span4Mux_v4 t1067 (
    .I(seg_13_12_sp4_v_b_9_50088),
    .O(seg_13_16_sp4_v_b_0_50573)
  );
  Span4Mux_v4 t1068 (
    .I(seg_13_8_sp4_v_b_9_49596),
    .O(seg_13_12_sp4_v_b_9_50088)
  );
  Span4Mux_v4 t1069 (
    .I(seg_13_4_sp4_h_l_44_37971),
    .O(seg_13_8_sp4_v_b_9_49596)
  );
  CascadeMux t107 (
    .I(net_38675),
    .O(net_38675_cascademuxed)
  );
  Span4Mux_h4 t1070 (
    .I(seg_9_4_sp4_v_b_3_33768),
    .O(seg_13_4_sp4_h_l_44_37971)
  );
  LocalMux t1071 (
    .I(seg_17_31_span4_vert_13_67863),
    .O(seg_17_31_local_g0_5_71851)
  );
  Span4Mux_v4 t1072 (
    .I(seg_17_28_sp4_v_b_9_67378),
    .O(seg_17_31_span4_vert_13_67863)
  );
  Span4Mux_v4 t1073 (
    .I(seg_17_24_sp4_v_b_6_66885),
    .O(seg_17_28_sp4_v_b_9_67378)
  );
  Span4Mux_v4 t1074 (
    .I(seg_17_20_sp4_v_b_6_66393),
    .O(seg_17_24_sp4_v_b_6_66885)
  );
  Span4Mux_v4 t1075 (
    .I(seg_17_16_sp4_v_b_6_65901),
    .O(seg_17_20_sp4_v_b_6_66393)
  );
  Span4Mux_v4 t1076 (
    .I(seg_17_12_sp4_v_b_3_65404),
    .O(seg_17_16_sp4_v_b_6_65901)
  );
  Span4Mux_v4 t1077 (
    .I(seg_17_8_sp4_v_b_0_64911),
    .O(seg_17_12_sp4_v_b_3_65404)
  );
  Span4Mux_v4 t1078 (
    .I(seg_17_4_sp4_h_l_37_53284),
    .O(seg_17_8_sp4_v_b_0_64911)
  );
  Span4Mux_h4 t1079 (
    .I(seg_13_4_sp4_h_l_44_37971),
    .O(seg_17_4_sp4_h_l_37_53284)
  );
  CascadeMux t108 (
    .I(net_38681),
    .O(net_38681_cascademuxed)
  );
  LocalMux t1080 (
    .I(seg_12_14_sp4_r_v_b_2_50329),
    .O(seg_12_14_local_g1_2_50599)
  );
  Span4Mux_v4 t1081 (
    .I(seg_13_10_sp4_v_b_11_49844),
    .O(seg_12_14_sp4_r_v_b_2_50329)
  );
  Span4Mux_v4 t1082 (
    .I(seg_13_6_sp4_h_l_46_38209),
    .O(seg_13_10_sp4_v_b_11_49844)
  );
  Span4Mux_h4 t1083 (
    .I(seg_9_6_sp4_v_b_11_34028),
    .O(seg_13_6_sp4_h_l_46_38209)
  );
  LocalMux t1084 (
    .I(seg_15_10_sp4_h_r_29_54029),
    .O(seg_15_10_local_g3_5_61617)
  );
  Span4Mux_h4 t1085 (
    .I(seg_13_10_sp4_v_b_11_49844),
    .O(seg_15_10_sp4_h_r_29_54029)
  );
  LocalMux t1086 (
    .I(seg_17_0_span4_vert_21_64396),
    .O(seg_17_0_local_g1_5_68058)
  );
  Span4Mux_v4 t1087 (
    .I(seg_17_2_sp4_h_l_39_53042),
    .O(seg_17_0_span4_vert_21_64396)
  );
  Span4Mux_h4 t1088 (
    .I(seg_13_2_sp4_h_l_46_37717),
    .O(seg_17_2_sp4_h_l_39_53042)
  );
  Span4Mux_h4 t1089 (
    .I(seg_9_2_sp4_v_t_46_34028),
    .O(seg_13_2_sp4_h_l_46_37717)
  );
  LocalMux t1090 (
    .I(seg_21_9_sp4_v_b_15_79852),
    .O(seg_21_9_local_g1_7_83835)
  );
  Span4Mux_v4 t1091 (
    .I(seg_21_6_sp4_h_l_39_68856),
    .O(seg_21_9_sp4_v_b_15_79852)
  );
  Span4Mux_h4 t1092 (
    .I(seg_17_6_sp4_h_l_46_53533),
    .O(seg_21_6_sp4_h_l_39_68856)
  );
  Span4Mux_h4 t1093 (
    .I(seg_13_6_sp4_h_l_46_38209),
    .O(seg_17_6_sp4_h_l_46_53533)
  );
  LocalMux t1094 (
    .I(seg_4_13_sp4_v_b_12_16478),
    .O(seg_4_13_local_g1_4_20461)
  );
  Span4Mux_v4 t1095 (
    .I(seg_4_10_sp4_h_r_1_20175),
    .O(seg_4_13_sp4_v_b_12_16478)
  );
  Span4Mux_h4 t1096 (
    .I(seg_8_10_sp4_v_b_1_30679),
    .O(seg_4_10_sp4_h_r_1_20175)
  );
  Span4Mux_v4 t1097 (
    .I(seg_8_6_sp4_v_b_10_30198),
    .O(seg_8_10_sp4_v_b_1_30679)
  );
  LocalMux t1098 (
    .I(seg_4_18_sp4_v_b_6_16977),
    .O(seg_4_18_local_g1_6_21078)
  );
  Span4Mux_v4 t1099 (
    .I(seg_4_14_sp4_h_r_6_20674),
    .O(seg_4_18_sp4_v_b_6_16977)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t110 (
    .carryinitin(),
    .carryinitout(t109)
  );
  Span4Mux_h4 t1100 (
    .I(seg_8_14_sp4_v_b_1_31171),
    .O(seg_4_14_sp4_h_r_6_20674)
  );
  Span4Mux_v4 t1101 (
    .I(seg_8_10_sp4_v_b_1_30679),
    .O(seg_8_14_sp4_v_b_1_31171)
  );
  LocalMux t1102 (
    .I(seg_11_17_sp4_r_v_b_13_46988),
    .O(seg_11_17_local_g2_5_47148)
  );
  Span4Mux_v4 t1103 (
    .I(seg_12_14_sp4_v_b_0_46496),
    .O(seg_11_17_sp4_r_v_b_13_46988)
  );
  Span4Mux_v4 t1104 (
    .I(seg_12_10_sp4_v_b_4_46008),
    .O(seg_12_14_sp4_v_b_0_46496)
  );
  Span4Mux_v4 t1105 (
    .I(seg_12_6_sp4_h_l_41_34381),
    .O(seg_12_10_sp4_v_b_4_46008)
  );
  Span4Mux_h4 t1106 (
    .I(seg_8_6_sp4_v_b_10_30198),
    .O(seg_12_6_sp4_h_l_41_34381)
  );
  LocalMux t1107 (
    .I(seg_19_13_sp4_r_v_b_19_76916),
    .O(seg_19_13_local_g3_3_77054)
  );
  Span4Mux_v4 t1108 (
    .I(seg_20_10_sp4_v_b_3_76503),
    .O(seg_19_13_sp4_r_v_b_19_76916)
  );
  Span4Mux_v4 t1109 (
    .I(seg_20_6_sp4_h_l_38_65026),
    .O(seg_20_10_sp4_v_b_3_76503)
  );
  CascadeMux t111 (
    .I(net_38891),
    .O(net_38891_cascademuxed)
  );
  Span4Mux_h4 t1110 (
    .I(seg_16_6_sp4_h_l_42_49708),
    .O(seg_20_6_sp4_h_l_38_65026)
  );
  Span4Mux_h4 t1111 (
    .I(seg_12_6_sp4_h_l_41_34381),
    .O(seg_16_6_sp4_h_l_42_49708)
  );
  LocalMux t1112 (
    .I(seg_19_13_sp4_r_v_b_21_76918),
    .O(seg_19_13_local_g3_5_77056)
  );
  Span4Mux_v4 t1113 (
    .I(seg_20_10_sp4_v_b_8_76510),
    .O(seg_19_13_sp4_r_v_b_21_76918)
  );
  Span4Mux_v4 t1114 (
    .I(seg_20_6_sp4_h_l_38_65026),
    .O(seg_20_10_sp4_v_b_8_76510)
  );
  LocalMux t1115 (
    .I(seg_19_14_sp4_r_v_b_5_76913),
    .O(seg_19_14_local_g1_5_77142)
  );
  Span4Mux_v4 t1116 (
    .I(seg_20_10_sp4_v_b_9_76509),
    .O(seg_19_14_sp4_r_v_b_5_76913)
  );
  Span4Mux_v4 t1117 (
    .I(seg_20_6_sp4_h_l_41_65027),
    .O(seg_20_10_sp4_v_b_9_76509)
  );
  Span4Mux_h4 t1118 (
    .I(seg_16_6_sp4_h_l_41_49705),
    .O(seg_20_6_sp4_h_l_41_65027)
  );
  Span4Mux_h4 t1119 (
    .I(seg_12_6_sp4_h_l_41_34381),
    .O(seg_16_6_sp4_h_l_41_49705)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t112 (
    .carryinitin(net_42755),
    .carryinitout(net_42799)
  );
  LocalMux t1120 (
    .I(seg_19_17_sp4_r_v_b_19_77324),
    .O(seg_19_17_local_g3_3_77462)
  );
  Span4Mux_v4 t1121 (
    .I(seg_20_14_sp4_v_b_6_76916),
    .O(seg_19_17_sp4_r_v_b_19_77324)
  );
  Span4Mux_v4 t1122 (
    .I(seg_20_10_sp4_v_b_3_76503),
    .O(seg_20_14_sp4_v_b_6_76916)
  );
  LocalMux t1123 (
    .I(seg_19_17_sp4_r_v_b_21_77326),
    .O(seg_19_17_local_g3_5_77464)
  );
  Span4Mux_v4 t1124 (
    .I(seg_20_14_sp4_v_b_8_76918),
    .O(seg_19_17_sp4_r_v_b_21_77326)
  );
  Span4Mux_v4 t1125 (
    .I(seg_20_10_sp4_v_b_8_76510),
    .O(seg_20_14_sp4_v_b_8_76918)
  );
  LocalMux t1126 (
    .I(seg_21_10_sp4_h_r_20_80217),
    .O(seg_21_10_local_g0_4_83947)
  );
  Span4Mux_h4 t1127 (
    .I(seg_20_10_sp4_v_b_3_76503),
    .O(seg_21_10_sp4_h_r_20_80217)
  );
  LocalMux t1128 (
    .I(seg_8_10_lutff_2_out_30903),
    .O(seg_8_10_local_g0_2_34775)
  );
  LocalMux t1129 (
    .I(seg_8_10_lutff_3_out_30904),
    .O(seg_8_10_local_g3_3_34800)
  );
  LocalMux t1130 (
    .I(seg_8_10_lutff_4_out_30905),
    .O(seg_8_10_local_g3_4_34801)
  );
  LocalMux t1131 (
    .I(seg_8_10_lutff_5_out_30906),
    .O(seg_8_10_local_g0_5_34778)
  );
  LocalMux t1132 (
    .I(seg_8_10_lutff_6_out_30907),
    .O(seg_8_10_local_g0_6_34779)
  );
  LocalMux t1133 (
    .I(seg_8_11_sp12_v_b_13_34250),
    .O(seg_8_11_local_g3_5_34925)
  );
  LocalMux t1134 (
    .I(seg_8_10_sp4_h_r_20_31047),
    .O(seg_8_10_local_g0_4_34777)
  );
  Span4Mux_h4 t1135 (
    .I(seg_7_10_sp4_v_b_3_27333),
    .O(seg_8_10_sp4_h_r_20_31047)
  );
  Span4Mux_v4 t1136 (
    .I(seg_7_10_sp4_h_r_3_31041),
    .O(seg_7_10_sp4_v_b_3_27333)
  );
  LocalMux t1137 (
    .I(seg_17_18_sp4_r_v_b_1_69971),
    .O(seg_17_18_local_g1_1_70243)
  );
  Span4Mux_v4 t1138 (
    .I(seg_18_14_sp4_v_b_5_69483),
    .O(seg_17_18_sp4_r_v_b_1_69971)
  );
  Span4Mux_v4 t1139 (
    .I(seg_18_10_sp4_h_l_40_57859),
    .O(seg_18_14_sp4_v_b_5_69483)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t114 (
    .carryinitin(),
    .carryinitout(t113)
  );
  Span4Mux_h4 t1140 (
    .I(seg_14_10_sp4_h_l_39_42533),
    .O(seg_18_10_sp4_h_l_40_57859)
  );
  Span4Mux_h4 t1141 (
    .I(seg_10_10_sp4_h_l_43_27633),
    .O(seg_14_10_sp4_h_l_39_42533)
  );
  LocalMux t1142 (
    .I(seg_8_12_sp4_r_v_b_28_35007),
    .O(seg_8_12_local_g0_4_35023)
  );
  Span4Mux_v4 t1143 (
    .I(seg_9_10_sp4_h_l_46_24008),
    .O(seg_8_12_sp4_r_v_b_28_35007)
  );
  LocalMux t1144 (
    .I(seg_8_10_neigh_op_top_5_31029),
    .O(seg_8_10_local_g1_5_34786)
  );
  LocalMux t1145 (
    .I(seg_8_11_lutff_5_out_31029),
    .O(seg_8_11_local_g0_5_34901)
  );
  LocalMux t1146 (
    .I(seg_8_12_lutff_1_out_31148),
    .O(seg_8_12_local_g0_1_35020)
  );
  LocalMux t1147 (
    .I(seg_8_11_sp4_v_b_18_30931),
    .O(seg_8_11_local_g0_2_34898)
  );
  Span4Mux_v4 t1148 (
    .I(seg_8_12_sp4_h_r_2_35117),
    .O(seg_8_11_sp4_v_b_18_30931)
  );
  LocalMux t1149 (
    .I(seg_8_10_sp4_v_b_26_30928),
    .O(seg_8_10_local_g3_2_34799)
  );
  LocalMux t1150 (
    .I(seg_9_29_sp4_r_v_b_1_40678),
    .O(seg_9_29_local_g1_1_40950)
  );
  Span4Mux_v4 t1151 (
    .I(seg_10_25_sp4_v_b_10_40197),
    .O(seg_9_29_sp4_r_v_b_1_40678)
  );
  Span4Mux_v4 t1152 (
    .I(seg_10_21_sp4_v_b_2_39697),
    .O(seg_10_25_sp4_v_b_10_40197)
  );
  Span4Mux_v4 t1153 (
    .I(seg_10_17_sp4_h_l_39_28343),
    .O(seg_10_21_sp4_v_b_2_39697)
  );
  LocalMux t1154 (
    .I(seg_10_26_sp4_v_b_43_40685),
    .O(seg_10_26_local_g3_3_44430)
  );
  Span4Mux_v4 t1155 (
    .I(seg_10_25_sp4_v_b_10_40197),
    .O(seg_10_26_sp4_v_b_43_40685)
  );
  LocalMux t1156 (
    .I(seg_10_29_sp4_v_b_1_40678),
    .O(seg_10_29_local_g0_1_44773)
  );
  Span4Mux_v4 t1157 (
    .I(seg_10_25_sp4_v_b_10_40197),
    .O(seg_10_29_sp4_v_b_1_40678)
  );
  LocalMux t1158 (
    .I(seg_9_28_sp4_v_b_2_36727),
    .O(seg_9_28_local_g1_2_40828)
  );
  Span4Mux_v4 t1159 (
    .I(seg_9_24_sp4_v_b_2_36235),
    .O(seg_9_28_sp4_v_b_2_36727)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t116 (
    .carryinitin(net_43370),
    .carryinitout(net_43414)
  );
  Span4Mux_v4 t1160 (
    .I(seg_9_20_sp4_v_b_6_35747),
    .O(seg_9_24_sp4_v_b_2_36235)
  );
  LocalMux t1161 (
    .I(seg_9_30_sp4_v_b_26_37219),
    .O(seg_9_30_local_g2_2_41082)
  );
  Span4Mux_v4 t1162 (
    .I(seg_9_28_sp4_v_b_2_36727),
    .O(seg_9_30_sp4_v_b_26_37219)
  );
  LocalMux t1163 (
    .I(seg_8_23_lutff_5_out_32505),
    .O(seg_8_23_local_g3_5_36401)
  );
  LocalMux t1164 (
    .I(seg_8_24_sp4_v_b_18_32530),
    .O(seg_8_24_local_g0_2_36497)
  );
  Span4Mux_v4 t1165 (
    .I(seg_8_25_sp4_h_r_2_36716),
    .O(seg_8_24_sp4_v_b_18_32530)
  );
  Span4Mux_h4 t1166 (
    .I(seg_8_25_sp4_v_b_2_32527),
    .O(seg_8_25_sp4_h_r_2_36716)
  );
  LocalMux t1167 (
    .I(seg_8_25_sp4_v_b_2_32527),
    .O(seg_8_25_local_g1_2_36628)
  );
  LocalMux t1168 (
    .I(seg_8_24_lutff_6_out_32629),
    .O(seg_8_24_local_g2_6_36517)
  );
  LocalMux t1169 (
    .I(seg_8_25_neigh_op_bot_6_32629),
    .O(seg_8_25_local_g0_6_36624)
  );
  CascadeMux t117 (
    .I(net_39629),
    .O(net_39629_cascademuxed)
  );
  LocalMux t1170 (
    .I(seg_8_25_lutff_2_out_32748),
    .O(seg_8_25_local_g2_2_36636)
  );
  LocalMux t1171 (
    .I(seg_8_25_lutff_3_out_32749),
    .O(seg_8_25_local_g0_3_36621)
  );
  LocalMux t1172 (
    .I(seg_8_25_lutff_4_out_32750),
    .O(seg_8_25_local_g1_4_36630)
  );
  LocalMux t1173 (
    .I(seg_8_25_lutff_5_out_32751),
    .O(seg_8_25_local_g3_5_36647)
  );
  LocalMux t1174 (
    .I(seg_8_25_lutff_7_out_32753),
    .O(seg_8_25_local_g1_7_36633)
  );
  LocalMux t1175 (
    .I(seg_8_25_sp4_h_r_12_32882),
    .O(seg_8_25_local_g0_4_36622)
  );
  LocalMux t1176 (
    .I(seg_12_23_sp4_h_r_47_40299),
    .O(seg_12_23_local_g2_7_51719)
  );
  Span4Mux_h4 t1177 (
    .I(seg_9_23_sp4_v_t_40_36605),
    .O(seg_12_23_sp4_h_r_47_40299)
  );
  LocalMux t1178 (
    .I(seg_8_23_sp4_h_r_4_36472),
    .O(seg_8_23_local_g0_4_36376)
  );
  Span4Mux_h4 t1179 (
    .I(seg_8_23_sp4_v_t_41_32775),
    .O(seg_8_23_sp4_h_r_4_36472)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t118 (
    .carryinitin(net_43493),
    .carryinitout(net_43537)
  );
  LocalMux t1180 (
    .I(seg_8_24_sp4_v_b_5_32405),
    .O(seg_8_24_local_g1_5_36508)
  );
  Span4Mux_v4 t1181 (
    .I(seg_8_24_sp4_v_t_44_32901),
    .O(seg_8_24_sp4_v_b_5_32405)
  );
  LocalMux t1182 (
    .I(seg_9_30_neigh_op_tnl_6_33486),
    .O(seg_9_30_local_g3_6_41094)
  );
  LocalMux t1183 (
    .I(seg_10_30_sp4_r_v_b_24_44879),
    .O(seg_10_30_local_g0_0_44895)
  );
  IoSpan4Mux t1184 (
    .I(seg_11_31_span4_horz_l_14_33556),
    .O(seg_10_30_sp4_r_v_b_24_44879)
  );
  LocalMux t1185 (
    .I(seg_10_30_sp4_h_r_30_37331),
    .O(seg_10_30_local_g3_6_44925)
  );
  Span4Mux_h4 t1186 (
    .I(seg_8_30_sp4_v_t_36_37347),
    .O(seg_10_30_sp4_h_r_30_37331)
  );
  LocalMux t1187 (
    .I(seg_8_2_neigh_op_rgt_0_33712),
    .O(seg_8_2_local_g2_0_33805)
  );
  LocalMux t1188 (
    .I(seg_9_2_lutff_1_out_33713),
    .O(seg_9_2_local_g2_1_37637)
  );
  LocalMux t1189 (
    .I(seg_9_2_lutff_2_out_33714),
    .O(seg_9_2_local_g2_2_37638)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t119 (
    .carryinitin(net_43616),
    .carryinitout(net_43660)
  );
  LocalMux t1190 (
    .I(seg_9_2_lutff_3_out_33715),
    .O(seg_9_2_local_g1_3_37631)
  );
  LocalMux t1191 (
    .I(seg_9_2_lutff_4_out_33716),
    .O(seg_9_2_local_g0_4_37624)
  );
  LocalMux t1192 (
    .I(seg_10_2_neigh_op_lft_4_33716),
    .O(seg_10_2_local_g0_4_41455)
  );
  LocalMux t1193 (
    .I(seg_10_3_neigh_op_bnl_4_33716),
    .O(seg_10_3_local_g2_4_41594)
  );
  LocalMux t1194 (
    .I(seg_9_2_lutff_5_out_33717),
    .O(seg_9_2_local_g1_5_37633)
  );
  LocalMux t1195 (
    .I(seg_9_3_neigh_op_bot_6_33718),
    .O(seg_9_3_local_g0_6_37749)
  );
  LocalMux t1196 (
    .I(seg_9_2_lutff_7_out_33719),
    .O(seg_9_2_local_g0_7_37627)
  );
  LocalMux t1197 (
    .I(seg_9_4_neigh_op_bot_0_33871),
    .O(seg_9_4_local_g0_0_37866)
  );
  LocalMux t1198 (
    .I(seg_8_2_neigh_op_tnr_1_33872),
    .O(seg_8_2_local_g3_1_33814)
  );
  LocalMux t1199 (
    .I(seg_8_3_neigh_op_rgt_1_33872),
    .O(seg_8_3_local_g2_1_33929)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t12 (
    .carryinitin(),
    .carryinitout(t11)
  );
  LocalMux t1200 (
    .I(seg_9_2_neigh_op_top_1_33872),
    .O(seg_9_2_local_g0_1_37621)
  );
  LocalMux t1201 (
    .I(seg_9_3_lutff_1_out_33872),
    .O(seg_9_3_local_g1_1_37752)
  );
  LocalMux t1202 (
    .I(seg_9_3_lutff_1_out_33872),
    .O(seg_9_3_local_g2_1_37760)
  );
  LocalMux t1203 (
    .I(seg_8_2_neigh_op_tnr_2_33873),
    .O(seg_8_2_local_g3_2_33815)
  );
  LocalMux t1204 (
    .I(seg_8_3_neigh_op_rgt_2_33873),
    .O(seg_8_3_local_g3_2_33938)
  );
  LocalMux t1205 (
    .I(seg_9_2_neigh_op_top_2_33873),
    .O(seg_9_2_local_g0_2_37622)
  );
  LocalMux t1206 (
    .I(seg_9_3_lutff_2_out_33873),
    .O(seg_9_3_local_g3_2_37769)
  );
  LocalMux t1207 (
    .I(seg_9_3_lutff_3_out_33874),
    .O(seg_9_3_local_g3_3_37770)
  );
  LocalMux t1208 (
    .I(seg_8_2_neigh_op_tnr_4_33875),
    .O(seg_8_2_local_g3_4_33817)
  );
  LocalMux t1209 (
    .I(seg_8_3_neigh_op_rgt_4_33875),
    .O(seg_8_3_local_g2_4_33932)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t121 (
    .carryinitin(),
    .carryinitout(t120)
  );
  LocalMux t1210 (
    .I(seg_9_2_neigh_op_top_4_33875),
    .O(seg_9_2_local_g1_4_37632)
  );
  LocalMux t1211 (
    .I(seg_9_3_lutff_4_out_33875),
    .O(seg_9_3_local_g1_4_37755)
  );
  LocalMux t1212 (
    .I(seg_9_3_lutff_4_out_33875),
    .O(seg_9_3_local_g2_4_37763)
  );
  LocalMux t1213 (
    .I(seg_9_3_lutff_5_out_33876),
    .O(seg_9_3_local_g2_5_37764)
  );
  LocalMux t1214 (
    .I(seg_9_3_lutff_6_out_33877),
    .O(seg_9_3_local_g1_6_37757)
  );
  LocalMux t1215 (
    .I(seg_9_2_neigh_op_top_7_33878),
    .O(seg_9_2_local_g1_7_37635)
  );
  LocalMux t1216 (
    .I(seg_9_3_lutff_7_out_33878),
    .O(seg_9_3_local_g2_7_37766)
  );
  LocalMux t1217 (
    .I(seg_9_4_lutff_1_out_33995),
    .O(seg_9_4_local_g2_1_37883)
  );
  LocalMux t1218 (
    .I(seg_9_3_neigh_op_top_5_33999),
    .O(seg_9_3_local_g1_5_37756)
  );
  LocalMux t1219 (
    .I(seg_9_5_sp4_h_r_11_38086),
    .O(seg_9_5_local_g1_3_38000)
  );
  Span4Mux_h4 t1220 (
    .I(seg_9_5_sp4_v_b_5_33899),
    .O(seg_9_5_sp4_h_r_11_38086)
  );
  LocalMux t1221 (
    .I(seg_9_10_sp4_r_v_b_10_38352),
    .O(seg_9_10_local_g2_2_38622)
  );
  Span4Mux_v4 t1222 (
    .I(seg_10_6_sp4_v_b_10_37860),
    .O(seg_9_10_sp4_r_v_b_10_38352)
  );
  LocalMux t1223 (
    .I(seg_10_10_sp4_v_b_6_38348),
    .O(seg_10_10_local_g0_6_42441)
  );
  Span4Mux_v4 t1224 (
    .I(seg_10_6_sp4_v_b_10_37860),
    .O(seg_10_10_sp4_v_b_6_38348)
  );
  LocalMux t1225 (
    .I(seg_11_10_sp4_h_r_13_42529),
    .O(seg_11_10_local_g0_5_46271)
  );
  Span4Mux_h4 t1226 (
    .I(seg_10_10_sp4_v_b_6_38348),
    .O(seg_11_10_sp4_h_r_13_42529)
  );
  LocalMux t1227 (
    .I(seg_10_8_neigh_op_lft_5_34491),
    .O(seg_10_8_local_g0_5_42194)
  );
  LocalMux t1228 (
    .I(seg_10_8_neigh_op_lft_6_34492),
    .O(seg_10_8_local_g1_6_42203)
  );
  LocalMux t1229 (
    .I(seg_10_8_neigh_op_lft_7_34493),
    .O(seg_10_8_local_g0_7_42196)
  );
  CascadeMux t123 (
    .I(net_40736),
    .O(net_40736_cascademuxed)
  );
  LocalMux t1230 (
    .I(seg_11_9_sp4_v_b_40_42422),
    .O(seg_11_9_local_g3_0_46167)
  );
  Span4Mux_v4 t1231 (
    .I(seg_11_8_sp4_h_l_37_30790),
    .O(seg_11_9_sp4_v_b_40_42422)
  );
  LocalMux t1232 (
    .I(seg_11_9_sp4_h_r_15_42410),
    .O(seg_11_9_local_g0_7_46150)
  );
  Span4Mux_h4 t1233 (
    .I(seg_10_9_sp4_v_b_8_38227),
    .O(seg_11_9_sp4_h_r_15_42410)
  );
  LocalMux t1234 (
    .I(seg_11_9_sp4_h_r_23_42408),
    .O(seg_11_9_local_g1_7_46158)
  );
  Span4Mux_h4 t1235 (
    .I(seg_10_9_sp4_v_b_10_38229),
    .O(seg_11_9_sp4_h_r_23_42408)
  );
  LocalMux t1236 (
    .I(seg_10_10_neigh_op_lft_1_34733),
    .O(seg_10_10_local_g0_1_42436)
  );
  LocalMux t1237 (
    .I(seg_9_10_lutff_2_out_34734),
    .O(seg_9_10_local_g3_2_38630)
  );
  LocalMux t1238 (
    .I(seg_9_10_lutff_4_out_34736),
    .O(seg_9_10_local_g3_4_38632)
  );
  LocalMux t1239 (
    .I(seg_10_11_neigh_op_bnl_4_34736),
    .O(seg_10_11_local_g3_4_42586)
  );
  CascadeMux t124 (
    .I(net_40760),
    .O(net_40760_cascademuxed)
  );
  LocalMux t1240 (
    .I(seg_9_10_lutff_7_out_34739),
    .O(seg_9_10_local_g2_7_38627)
  );
  LocalMux t1241 (
    .I(seg_11_10_sp4_h_r_36_34868),
    .O(seg_11_10_local_g2_4_46286)
  );
  LocalMux t1242 (
    .I(seg_11_10_sp4_h_r_36_34868),
    .O(seg_11_10_local_g3_4_46294)
  );
  LocalMux t1243 (
    .I(seg_11_10_sp4_h_r_26_38702),
    .O(seg_11_10_local_g3_2_46292)
  );
  LocalMux t1244 (
    .I(seg_10_12_sp4_v_b_17_38715),
    .O(seg_10_12_local_g1_1_42690)
  );
  LocalMux t1245 (
    .I(seg_10_11_neigh_op_lft_5_34860),
    .O(seg_10_11_local_g0_5_42563)
  );
  LocalMux t1246 (
    .I(seg_13_14_sp4_v_b_23_50460),
    .O(seg_13_14_local_g1_7_54435)
  );
  Span4Mux_v4 t1247 (
    .I(seg_13_11_sp4_h_l_47_38823),
    .O(seg_13_14_sp4_v_b_23_50460)
  );
  LocalMux t1248 (
    .I(seg_13_3_sp4_r_v_b_23_52933),
    .O(seg_13_3_local_g3_7_53098)
  );
  Span4Mux_v4 t1249 (
    .I(seg_14_4_sp4_h_l_41_41797),
    .O(seg_13_3_sp4_r_v_b_23_52933)
  );
  CascadeMux t125 (
    .I(net_40859),
    .O(net_40859_cascademuxed)
  );
  Span4Mux_h4 t1250 (
    .I(seg_10_4_sp4_v_t_46_38105),
    .O(seg_14_4_sp4_h_l_41_41797)
  );
  Span4Mux_v4 t1251 (
    .I(seg_10_8_sp4_v_t_38_38589),
    .O(seg_10_4_sp4_v_t_46_38105)
  );
  LocalMux t1252 (
    .I(seg_14_3_sp4_v_b_14_52923),
    .O(seg_14_3_local_g1_6_56911)
  );
  Span4Mux_v4 t1253 (
    .I(seg_14_4_sp4_v_t_38_53421),
    .O(seg_14_3_sp4_v_b_14_52923)
  );
  Span4Mux_v4 t1254 (
    .I(seg_14_8_sp4_h_l_38_42288),
    .O(seg_14_4_sp4_v_t_38_53421)
  );
  Span4Mux_h4 t1255 (
    .I(seg_10_8_sp4_v_t_38_38589),
    .O(seg_14_8_sp4_h_l_38_42288)
  );
  LocalMux t1256 (
    .I(seg_10_26_sp4_v_b_10_40320),
    .O(seg_10_26_local_g1_2_44413)
  );
  Span4Mux_v4 t1257 (
    .I(seg_10_22_sp4_v_b_10_39828),
    .O(seg_10_26_sp4_v_b_10_40320)
  );
  Span4Mux_v4 t1258 (
    .I(seg_10_18_sp4_v_b_7_39331),
    .O(seg_10_22_sp4_v_b_10_39828)
  );
  Span4Mux_v4 t1259 (
    .I(seg_10_14_sp4_v_b_11_38843),
    .O(seg_10_18_sp4_v_b_7_39331)
  );
  CascadeMux t126 (
    .I(net_40865),
    .O(net_40865_cascademuxed)
  );
  LocalMux t1260 (
    .I(seg_14_26_sp4_v_b_9_55641),
    .O(seg_14_26_local_g1_1_59735)
  );
  Span4Mux_v4 t1261 (
    .I(seg_14_22_sp4_v_b_6_55148),
    .O(seg_14_26_sp4_v_b_9_55641)
  );
  Span4Mux_v4 t1262 (
    .I(seg_14_18_sp4_v_b_10_54660),
    .O(seg_14_22_sp4_v_b_6_55148)
  );
  Span4Mux_v4 t1263 (
    .I(seg_14_14_sp4_h_l_40_43028),
    .O(seg_14_18_sp4_v_b_10_54660)
  );
  Span4Mux_h4 t1264 (
    .I(seg_10_14_sp4_v_b_11_38843),
    .O(seg_14_14_sp4_h_l_40_43028)
  );
  LocalMux t1265 (
    .I(seg_9_4_sp4_h_r_3_37965),
    .O(seg_9_4_local_g0_3_37869)
  );
  Span4Mux_h4 t1266 (
    .I(seg_9_4_sp4_v_t_47_34275),
    .O(seg_9_4_sp4_h_r_3_37965)
  );
  Span4Mux_v4 t1267 (
    .I(seg_9_8_sp4_v_t_39_34759),
    .O(seg_9_4_sp4_v_t_47_34275)
  );
  LocalMux t1268 (
    .I(seg_11_18_sp4_h_r_26_39686),
    .O(seg_11_18_local_g3_2_47276)
  );
  LocalMux t1269 (
    .I(seg_11_18_sp4_h_r_16_43520),
    .O(seg_11_18_local_g1_0_47258)
  );
  CascadeMux t127 (
    .I(net_40889),
    .O(net_40889_cascademuxed)
  );
  Span4Mux_h4 t1270 (
    .I(seg_10_18_sp4_v_b_11_39335),
    .O(seg_11_18_sp4_h_r_16_43520)
  );
  LocalMux t1271 (
    .I(seg_9_27_lutff_1_out_36824),
    .O(seg_9_27_local_g0_1_40696)
  );
  LocalMux t1272 (
    .I(seg_9_28_neigh_op_bot_5_36828),
    .O(seg_9_28_local_g1_5_40831)
  );
  LocalMux t1273 (
    .I(seg_10_27_neigh_op_lft_5_36828),
    .O(seg_10_27_local_g0_5_44531)
  );
  LocalMux t1274 (
    .I(seg_10_28_neigh_op_bnl_5_36828),
    .O(seg_10_28_local_g2_5_44670)
  );
  LocalMux t1275 (
    .I(seg_9_27_lutff_7_out_36830),
    .O(seg_9_27_local_g2_7_40718)
  );
  LocalMux t1276 (
    .I(seg_9_28_neigh_op_bot_7_36830),
    .O(seg_9_28_local_g1_7_40833)
  );
  LocalMux t1277 (
    .I(seg_10_27_neigh_op_lft_7_36830),
    .O(seg_10_27_local_g1_7_44541)
  );
  LocalMux t1278 (
    .I(seg_10_28_neigh_op_bnl_7_36830),
    .O(seg_10_28_local_g3_7_44680)
  );
  LocalMux t1279 (
    .I(seg_9_28_lutff_2_out_36948),
    .O(seg_9_28_local_g0_2_40820)
  );
  CascadeMux t128 (
    .I(net_40976),
    .O(net_40976_cascademuxed)
  );
  LocalMux t1280 (
    .I(seg_9_28_lutff_5_out_36951),
    .O(seg_9_28_local_g2_5_40839)
  );
  LocalMux t1281 (
    .I(seg_9_28_sp4_h_r_34_33252),
    .O(seg_9_28_local_g2_2_40836)
  );
  LocalMux t1282 (
    .I(seg_9_30_sp4_v_b_20_37101),
    .O(seg_9_30_local_g0_4_41068)
  );
  LocalMux t1283 (
    .I(seg_9_29_lutff_0_out_37069),
    .O(seg_9_29_local_g0_0_40941)
  );
  LocalMux t1284 (
    .I(seg_10_28_neigh_op_tnl_3_37072),
    .O(seg_10_28_local_g3_3_44676)
  );
  LocalMux t1285 (
    .I(seg_9_28_neigh_op_top_5_37074),
    .O(seg_9_28_local_g0_5_40823)
  );
  LocalMux t1286 (
    .I(seg_9_27_sp4_r_v_b_27_40680),
    .O(seg_9_27_local_g1_3_40706)
  );
  Span4Mux_v4 t1287 (
    .I(seg_10_29_sp4_h_l_38_29568),
    .O(seg_9_27_sp4_r_v_b_27_40680)
  );
  LocalMux t1288 (
    .I(seg_10_27_sp4_v_b_27_40680),
    .O(seg_10_27_local_g3_3_44553)
  );
  Span4Mux_v4 t1289 (
    .I(seg_10_29_sp4_h_l_38_29568),
    .O(seg_10_27_sp4_v_b_27_40680)
  );
  CascadeMux t129 (
    .I(net_41006),
    .O(net_41006_cascademuxed)
  );
  LocalMux t1290 (
    .I(seg_9_30_lutff_0_out_37192),
    .O(seg_9_30_local_g0_0_41064)
  );
  LocalMux t1291 (
    .I(seg_10_30_neigh_op_lft_5_37197),
    .O(seg_10_30_local_g0_5_44900)
  );
  LocalMux t1292 (
    .I(seg_8_31_logic_op_bnr_7_37199),
    .O(seg_8_31_local_g0_7_37376)
  );
  LocalMux t1293 (
    .I(seg_10_2_lutff_2_out_37545),
    .O(seg_10_2_local_g3_2_41477)
  );
  LocalMux t1294 (
    .I(seg_10_3_neigh_op_bot_3_37546),
    .O(seg_10_3_local_g1_3_41585)
  );
  LocalMux t1295 (
    .I(seg_10_2_lutff_4_out_37547),
    .O(seg_10_2_local_g2_4_41471)
  );
  LocalMux t1296 (
    .I(seg_10_3_neigh_op_bot_5_37548),
    .O(seg_10_3_local_g1_5_41587)
  );
  LocalMux t1297 (
    .I(seg_9_2_neigh_op_rgt_6_37549),
    .O(seg_9_2_local_g3_6_37650)
  );
  LocalMux t1298 (
    .I(seg_10_2_lutff_6_out_37549),
    .O(seg_10_2_local_g1_6_41465)
  );
  LocalMux t1299 (
    .I(seg_9_2_neigh_op_rgt_7_37550),
    .O(seg_9_2_local_g2_7_37643)
  );
  CascadeMux t130 (
    .I(net_41099),
    .O(net_41099_cascademuxed)
  );
  LocalMux t1300 (
    .I(seg_9_2_neigh_op_rgt_7_37550),
    .O(seg_9_2_local_g3_7_37651)
  );
  LocalMux t1301 (
    .I(seg_10_2_lutff_7_out_37550),
    .O(seg_10_2_local_g0_7_41458)
  );
  LocalMux t1302 (
    .I(seg_9_2_neigh_op_tnr_2_37704),
    .O(seg_9_2_local_g3_2_37646)
  );
  LocalMux t1303 (
    .I(seg_10_2_neigh_op_top_2_37704),
    .O(seg_10_2_local_g0_2_41453)
  );
  LocalMux t1304 (
    .I(seg_9_2_neigh_op_tnr_3_37705),
    .O(seg_9_2_local_g3_3_37647)
  );
  LocalMux t1305 (
    .I(seg_10_2_neigh_op_top_3_37705),
    .O(seg_10_2_local_g0_3_41454)
  );
  LocalMux t1306 (
    .I(seg_10_3_lutff_3_out_37705),
    .O(seg_10_3_local_g3_3_41601)
  );
  LocalMux t1307 (
    .I(seg_9_2_neigh_op_tnr_4_37706),
    .O(seg_9_2_local_g2_4_37640)
  );
  LocalMux t1308 (
    .I(seg_10_2_neigh_op_top_4_37706),
    .O(seg_10_2_local_g1_4_41463)
  );
  LocalMux t1309 (
    .I(seg_9_2_neigh_op_tnr_6_37708),
    .O(seg_9_2_local_g2_6_37642)
  );
  CascadeMux t131 (
    .I(net_41111),
    .O(net_41111_cascademuxed)
  );
  LocalMux t1310 (
    .I(seg_10_2_neigh_op_top_6_37708),
    .O(seg_10_2_local_g0_6_41457)
  );
  LocalMux t1311 (
    .I(seg_10_3_lutff_6_out_37708),
    .O(seg_10_3_local_g1_6_41588)
  );
  LocalMux t1312 (
    .I(seg_10_3_lutff_7_out_37709),
    .O(seg_10_3_local_g3_7_41605)
  );
  LocalMux t1313 (
    .I(seg_14_7_sp4_h_r_10_57485),
    .O(seg_14_7_local_g0_2_57391)
  );
  Span4Mux_h4 t1314 (
    .I(seg_14_7_sp4_h_l_47_42162),
    .O(seg_14_7_sp4_h_r_10_57485)
  );
  LocalMux t1315 (
    .I(seg_14_8_sp4_v_b_43_53795),
    .O(seg_14_8_local_g3_3_57539)
  );
  Span4Mux_v4 t1316 (
    .I(seg_14_7_sp4_h_r_6_57491),
    .O(seg_14_8_sp4_v_b_43_53795)
  );
  Span4Mux_h4 t1317 (
    .I(seg_14_7_sp4_h_l_47_42162),
    .O(seg_14_7_sp4_h_r_6_57491)
  );
  LocalMux t1318 (
    .I(seg_11_7_sp4_v_b_11_41813),
    .O(seg_11_7_local_g1_3_45908)
  );
  LocalMux t1319 (
    .I(seg_11_9_sp4_v_b_3_42051),
    .O(seg_11_9_local_g1_3_46154)
  );
  CascadeMux t132 (
    .I(net_41504),
    .O(net_41504_cascademuxed)
  );
  LocalMux t1320 (
    .I(seg_13_9_sp4_h_r_27_46242),
    .O(seg_13_9_local_g3_3_53832)
  );
  Span4Mux_h4 t1321 (
    .I(seg_11_9_sp4_v_b_3_42051),
    .O(seg_13_9_sp4_h_r_27_46242)
  );
  LocalMux t1322 (
    .I(seg_10_8_sp4_v_b_43_38471),
    .O(seg_10_8_local_g3_3_42216)
  );
  Span4Mux_v4 t1323 (
    .I(seg_10_7_sp4_v_b_10_37983),
    .O(seg_10_8_sp4_v_b_43_38471)
  );
  LocalMux t1324 (
    .I(seg_10_8_lutff_0_out_38317),
    .O(seg_10_8_local_g2_0_42205)
  );
  LocalMux t1325 (
    .I(seg_9_8_neigh_op_rgt_2_38319),
    .O(seg_9_8_local_g2_2_38376)
  );
  LocalMux t1326 (
    .I(seg_11_8_neigh_op_lft_2_38319),
    .O(seg_11_8_local_g0_2_46022)
  );
  LocalMux t1327 (
    .I(seg_10_8_lutff_3_out_38320),
    .O(seg_10_8_local_g1_3_42200)
  );
  LocalMux t1328 (
    .I(seg_9_8_neigh_op_rgt_4_38321),
    .O(seg_9_8_local_g3_4_38386)
  );
  LocalMux t1329 (
    .I(seg_11_8_neigh_op_lft_4_38321),
    .O(seg_11_8_local_g0_4_46024)
  );
  CascadeMux t133 (
    .I(net_41522),
    .O(net_41522_cascademuxed)
  );
  LocalMux t1330 (
    .I(seg_9_8_neigh_op_rgt_6_38323),
    .O(seg_9_8_local_g2_6_38380)
  );
  LocalMux t1331 (
    .I(seg_11_8_neigh_op_lft_6_38323),
    .O(seg_11_8_local_g1_6_46034)
  );
  LocalMux t1332 (
    .I(seg_10_8_lutff_7_out_38324),
    .O(seg_10_8_local_g2_7_42212)
  );
  LocalMux t1333 (
    .I(seg_11_10_sp4_v_b_11_42182),
    .O(seg_11_10_local_g1_3_46277)
  );
  LocalMux t1334 (
    .I(seg_10_11_neigh_op_bot_2_38565),
    .O(seg_10_11_local_g0_2_42560)
  );
  LocalMux t1335 (
    .I(seg_10_13_sp4_r_v_b_19_42671),
    .O(seg_10_13_local_g3_3_42831)
  );
  Span4Mux_v4 t1336 (
    .I(seg_11_10_sp4_h_l_36_31037),
    .O(seg_10_13_sp4_r_v_b_19_42671)
  );
  LocalMux t1337 (
    .I(seg_10_12_sp4_v_b_34_38844),
    .O(seg_10_12_local_g2_2_42699)
  );
  Span4Mux_v4 t1338 (
    .I(seg_10_10_sp4_h_r_4_42535),
    .O(seg_10_12_sp4_v_b_34_38844)
  );
  LocalMux t1339 (
    .I(seg_10_12_neigh_op_bot_0_38686),
    .O(seg_10_12_local_g1_0_42689)
  );
  CascadeMux t134 (
    .I(net_41621),
    .O(net_41621_cascademuxed)
  );
  LocalMux t1340 (
    .I(seg_10_12_neigh_op_bot_1_38687),
    .O(seg_10_12_local_g0_1_42682)
  );
  LocalMux t1341 (
    .I(seg_10_11_lutff_4_out_38690),
    .O(seg_10_11_local_g2_4_42578)
  );
  LocalMux t1342 (
    .I(seg_10_12_neigh_op_bot_4_38690),
    .O(seg_10_12_local_g1_4_42693)
  );
  LocalMux t1343 (
    .I(seg_12_14_sp4_h_r_19_46860),
    .O(seg_12_14_local_g1_3_50600)
  );
  Span4Mux_h4 t1344 (
    .I(seg_11_14_sp4_v_b_0_42665),
    .O(seg_12_14_sp4_h_r_19_46860)
  );
  LocalMux t1345 (
    .I(seg_11_12_neigh_op_lft_1_38810),
    .O(seg_11_12_local_g0_1_46513)
  );
  LocalMux t1346 (
    .I(seg_11_12_neigh_op_lft_5_38814),
    .O(seg_11_12_local_g0_5_46517)
  );
  LocalMux t1347 (
    .I(seg_11_12_neigh_op_lft_7_38816),
    .O(seg_11_12_local_g0_7_46519)
  );
  LocalMux t1348 (
    .I(seg_13_12_sp4_h_r_1_54269),
    .O(seg_13_12_local_g0_1_54175)
  );
  Span4Mux_h4 t1349 (
    .I(seg_13_12_sp4_h_l_36_38945),
    .O(seg_13_12_sp4_h_r_1_54269)
  );
  CascadeMux t135 (
    .I(net_41633),
    .O(net_41633_cascademuxed)
  );
  LocalMux t1350 (
    .I(seg_13_12_sp4_h_r_41_42781),
    .O(seg_13_12_local_g2_1_54191)
  );
  LocalMux t1351 (
    .I(seg_13_12_sp4_h_r_43_42783),
    .O(seg_13_12_local_g2_3_54193)
  );
  LocalMux t1352 (
    .I(seg_13_12_sp4_h_r_45_42785),
    .O(seg_13_12_local_g2_5_54195)
  );
  LocalMux t1353 (
    .I(seg_11_13_neigh_op_lft_1_38933),
    .O(seg_11_13_local_g1_1_46644)
  );
  LocalMux t1354 (
    .I(seg_11_13_neigh_op_lft_2_38934),
    .O(seg_11_13_local_g1_2_46645)
  );
  LocalMux t1355 (
    .I(seg_11_13_neigh_op_lft_4_38936),
    .O(seg_11_13_local_g0_4_46639)
  );
  LocalMux t1356 (
    .I(seg_11_13_neigh_op_lft_5_38937),
    .O(seg_11_13_local_g1_5_46648)
  );
  LocalMux t1357 (
    .I(seg_11_13_neigh_op_lft_6_38938),
    .O(seg_11_13_local_g0_6_46641)
  );
  LocalMux t1358 (
    .I(seg_11_13_neigh_op_lft_7_38939),
    .O(seg_11_13_local_g1_7_46650)
  );
  LocalMux t1359 (
    .I(seg_13_13_sp4_h_r_37_42898),
    .O(seg_13_13_local_g3_5_54326)
  );
  CascadeMux t136 (
    .I(net_41645),
    .O(net_41645_cascademuxed)
  );
  LocalMux t1360 (
    .I(seg_13_13_sp4_h_r_43_42906),
    .O(seg_13_13_local_g2_3_54316)
  );
  LocalMux t1361 (
    .I(seg_10_13_neigh_op_top_0_39055),
    .O(seg_10_13_local_g1_0_42812)
  );
  LocalMux t1362 (
    .I(seg_10_13_neigh_op_top_1_39056),
    .O(seg_10_13_local_g0_1_42805)
  );
  LocalMux t1363 (
    .I(seg_10_14_lutff_2_out_39057),
    .O(seg_10_14_local_g2_2_42945)
  );
  LocalMux t1364 (
    .I(seg_10_13_neigh_op_top_3_39058),
    .O(seg_10_13_local_g0_3_42807)
  );
  LocalMux t1365 (
    .I(seg_10_14_lutff_4_out_39059),
    .O(seg_10_14_local_g2_4_42947)
  );
  LocalMux t1366 (
    .I(seg_11_14_neigh_op_lft_4_39059),
    .O(seg_11_14_local_g0_4_46762)
  );
  LocalMux t1367 (
    .I(seg_10_14_lutff_6_out_39061),
    .O(seg_10_14_local_g1_6_42941)
  );
  LocalMux t1368 (
    .I(seg_11_14_neigh_op_lft_6_39061),
    .O(seg_11_14_local_g0_6_46764)
  );
  LocalMux t1369 (
    .I(seg_10_14_lutff_7_out_39062),
    .O(seg_10_14_local_g3_7_42958)
  );
  CascadeMux t137 (
    .I(net_41651),
    .O(net_41651_cascademuxed)
  );
  LocalMux t1370 (
    .I(seg_11_14_neigh_op_lft_7_39062),
    .O(seg_11_14_local_g1_7_46773)
  );
  LocalMux t1371 (
    .I(seg_12_14_sp4_h_r_28_43027),
    .O(seg_12_14_local_g2_4_50609)
  );
  LocalMux t1372 (
    .I(seg_10_12_sp4_r_v_b_35_42674),
    .O(seg_10_12_local_g2_3_42700)
  );
  LocalMux t1373 (
    .I(seg_10_15_lutff_2_out_39180),
    .O(seg_10_15_local_g0_2_43052)
  );
  LocalMux t1374 (
    .I(seg_12_15_sp4_h_r_28_43150),
    .O(seg_12_15_local_g3_4_50740)
  );
  LocalMux t1375 (
    .I(seg_10_13_sp4_v_b_24_38957),
    .O(seg_10_13_local_g3_0_42828)
  );
  LocalMux t1376 (
    .I(seg_10_12_sp4_v_b_45_38965),
    .O(seg_10_12_local_g2_5_42702)
  );
  LocalMux t1377 (
    .I(seg_10_17_lutff_2_out_39426),
    .O(seg_10_17_local_g3_2_43322)
  );
  LocalMux t1378 (
    .I(seg_10_17_lutff_3_out_39427),
    .O(seg_10_17_local_g2_3_43315)
  );
  LocalMux t1379 (
    .I(seg_10_17_lutff_4_out_39428),
    .O(seg_10_17_local_g0_4_43300)
  );
  LocalMux t1380 (
    .I(seg_10_17_lutff_5_out_39429),
    .O(seg_10_17_local_g3_5_43325)
  );
  LocalMux t1381 (
    .I(seg_10_17_lutff_6_out_39430),
    .O(seg_10_17_local_g0_6_43302)
  );
  LocalMux t1382 (
    .I(seg_10_17_lutff_7_out_39431),
    .O(seg_10_17_local_g1_7_43311)
  );
  LocalMux t1383 (
    .I(seg_12_13_sp4_r_v_b_9_50211),
    .O(seg_12_13_local_g2_1_50483)
  );
  Span4Mux_v4 t1384 (
    .I(seg_13_13_sp4_v_t_44_50703),
    .O(seg_12_13_sp4_r_v_b_9_50211)
  );
  Span4Mux_v4 t1385 (
    .I(seg_13_17_sp4_h_l_38_39564),
    .O(seg_13_13_sp4_v_t_44_50703)
  );
  LocalMux t1386 (
    .I(seg_12_17_sp4_h_r_38_39564),
    .O(seg_12_17_local_g2_6_50980)
  );
  LocalMux t1387 (
    .I(seg_13_17_sp4_h_r_6_54891),
    .O(seg_13_17_local_g1_6_54803)
  );
  Span4Mux_h4 t1388 (
    .I(seg_13_17_sp4_h_l_38_39564),
    .O(seg_13_17_sp4_h_r_6_54891)
  );
  LocalMux t1389 (
    .I(seg_16_15_sp4_r_v_b_24_66018),
    .O(seg_16_15_local_g0_0_66034)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t139 (
    .carryinitin(),
    .carryinitout(t138)
  );
  Span4Mux_v4 t1390 (
    .I(seg_17_17_sp4_h_l_37_54883),
    .O(seg_16_15_sp4_r_v_b_24_66018)
  );
  Span4Mux_h4 t1391 (
    .I(seg_13_17_sp4_h_l_44_39570),
    .O(seg_17_17_sp4_h_l_37_54883)
  );
  LocalMux t1392 (
    .I(seg_16_16_sp4_r_v_b_13_66018),
    .O(seg_16_16_local_g2_5_66178)
  );
  Span4Mux_v4 t1393 (
    .I(seg_17_17_sp4_h_l_37_54883),
    .O(seg_16_16_sp4_r_v_b_13_66018)
  );
  LocalMux t1394 (
    .I(seg_12_12_sp4_v_b_16_46376),
    .O(seg_12_12_local_g0_0_50343)
  );
  Span4Mux_v4 t1395 (
    .I(seg_12_13_sp4_v_t_39_46867),
    .O(seg_12_12_sp4_v_b_16_46376)
  );
  Span4Mux_v4 t1396 (
    .I(seg_12_17_sp4_h_l_39_35732),
    .O(seg_12_13_sp4_v_t_39_46867)
  );
  LocalMux t1397 (
    .I(seg_12_12_sp4_v_b_13_46373),
    .O(seg_12_12_local_g1_5_50356)
  );
  Span4Mux_v4 t1398 (
    .I(seg_12_13_sp4_v_t_41_46869),
    .O(seg_12_12_sp4_v_b_13_46373)
  );
  Span4Mux_v4 t1399 (
    .I(seg_12_17_sp4_h_l_41_35734),
    .O(seg_12_13_sp4_v_t_41_46869)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t14 (
    .carryinitin(net_17307),
    .carryinitout(net_17351)
  );
  LocalMux t1400 (
    .I(seg_16_12_sp4_v_b_15_61697),
    .O(seg_16_12_local_g1_7_65680)
  );
  Span4Mux_v4 t1401 (
    .I(seg_16_13_sp4_v_t_43_62193),
    .O(seg_16_12_sp4_v_b_15_61697)
  );
  Span4Mux_v4 t1402 (
    .I(seg_16_17_sp4_h_l_37_51052),
    .O(seg_16_13_sp4_v_t_43_62193)
  );
  Span4Mux_h4 t1403 (
    .I(seg_12_17_sp4_h_l_41_35734),
    .O(seg_16_17_sp4_h_l_37_51052)
  );
  LocalMux t1404 (
    .I(seg_14_11_sp4_v_b_30_54041),
    .O(seg_14_11_local_g2_6_57903)
  );
  Span4Mux_v4 t1405 (
    .I(seg_14_13_sp4_v_t_43_54533),
    .O(seg_14_11_sp4_v_b_30_54041)
  );
  Span4Mux_v4 t1406 (
    .I(seg_14_17_sp4_h_l_43_43398),
    .O(seg_14_13_sp4_v_t_43_54533)
  );
  LocalMux t1407 (
    .I(seg_14_12_sp4_v_b_19_54041),
    .O(seg_14_12_local_g0_3_58007)
  );
  Span4Mux_v4 t1408 (
    .I(seg_14_13_sp4_v_t_43_54533),
    .O(seg_14_12_sp4_v_b_19_54041)
  );
  LocalMux t1409 (
    .I(seg_14_15_sp4_v_b_30_54533),
    .O(seg_14_15_local_g2_6_58395)
  );
  CascadeMux t141 (
    .I(net_42224),
    .O(net_42224_cascademuxed)
  );
  Span4Mux_v4 t1410 (
    .I(seg_14_17_sp4_h_l_43_43398),
    .O(seg_14_15_sp4_v_b_30_54533)
  );
  LocalMux t1411 (
    .I(seg_13_16_sp4_r_v_b_21_54535),
    .O(seg_13_16_local_g3_5_54695)
  );
  Span4Mux_v4 t1412 (
    .I(seg_14_17_sp4_h_l_45_43400),
    .O(seg_13_16_sp4_r_v_b_21_54535)
  );
  LocalMux t1413 (
    .I(seg_11_11_sp4_v_b_26_42544),
    .O(seg_11_11_local_g2_2_46407)
  );
  Span4Mux_v4 t1414 (
    .I(seg_11_13_sp4_v_t_46_43043),
    .O(seg_11_11_sp4_v_b_26_42544)
  );
  LocalMux t1415 (
    .I(seg_14_11_sp4_r_v_b_35_57874),
    .O(seg_14_11_local_g2_3_57900)
  );
  Span4Mux_v4 t1416 (
    .I(seg_15_13_sp4_h_l_46_46732),
    .O(seg_14_11_sp4_r_v_b_35_57874)
  );
  Span4Mux_h4 t1417 (
    .I(seg_11_13_sp4_v_t_46_43043),
    .O(seg_15_13_sp4_h_l_46_46732)
  );
  LocalMux t1418 (
    .I(seg_15_11_sp4_v_b_35_57874),
    .O(seg_15_11_local_g2_3_61730)
  );
  Span4Mux_v4 t1419 (
    .I(seg_15_13_sp4_h_l_46_46732),
    .O(seg_15_11_sp4_v_b_35_57874)
  );
  CascadeMux t142 (
    .I(net_42230),
    .O(net_42230_cascademuxed)
  );
  LocalMux t1420 (
    .I(seg_14_12_sp4_r_v_b_30_57994),
    .O(seg_14_12_local_g1_6_58018)
  );
  Span4Mux_v4 t1421 (
    .I(seg_15_14_sp4_h_l_37_46852),
    .O(seg_14_12_sp4_r_v_b_30_57994)
  );
  Span4Mux_h4 t1422 (
    .I(seg_11_14_sp4_v_t_37_43157),
    .O(seg_15_14_sp4_h_l_37_46852)
  );
  LocalMux t1423 (
    .I(seg_15_11_sp4_v_b_43_57994),
    .O(seg_15_11_local_g3_3_61738)
  );
  Span4Mux_v4 t1424 (
    .I(seg_15_14_sp4_h_l_37_46852),
    .O(seg_15_11_sp4_v_b_43_57994)
  );
  LocalMux t1425 (
    .I(seg_16_14_sp4_h_r_14_62179),
    .O(seg_16_14_local_g0_6_65917)
  );
  Span4Mux_h4 t1426 (
    .I(seg_15_14_sp4_h_l_37_46852),
    .O(seg_16_14_sp4_h_r_14_62179)
  );
  LocalMux t1427 (
    .I(seg_11_14_sp4_h_r_7_46861),
    .O(seg_11_14_local_g0_7_46765)
  );
  Span4Mux_h4 t1428 (
    .I(seg_11_14_sp4_v_t_39_43159),
    .O(seg_11_14_sp4_h_r_7_46861)
  );
  LocalMux t1429 (
    .I(seg_15_15_sp4_h_r_6_62305),
    .O(seg_15_15_local_g1_6_62217)
  );
  CascadeMux t143 (
    .I(net_42242),
    .O(net_42242_cascademuxed)
  );
  Span4Mux_h4 t1430 (
    .I(seg_15_15_sp4_h_l_43_46983),
    .O(seg_15_15_sp4_h_r_6_62305)
  );
  Span4Mux_h4 t1431 (
    .I(seg_11_15_sp4_v_t_36_43279),
    .O(seg_15_15_sp4_h_l_43_46983)
  );
  LocalMux t1432 (
    .I(seg_12_11_sp4_h_r_17_46489),
    .O(seg_12_11_local_g1_1_50229)
  );
  Span4Mux_h4 t1433 (
    .I(seg_11_11_sp4_v_t_46_42797),
    .O(seg_12_11_sp4_h_r_17_46489)
  );
  Span4Mux_v4 t1434 (
    .I(seg_11_15_sp4_v_t_38_43281),
    .O(seg_11_11_sp4_v_t_46_42797)
  );
  LocalMux t1435 (
    .I(seg_14_15_sp4_h_r_45_46985),
    .O(seg_14_15_local_g3_5_58402)
  );
  Span4Mux_h4 t1436 (
    .I(seg_11_15_sp4_v_t_38_43281),
    .O(seg_14_15_sp4_h_r_45_46985)
  );
  LocalMux t1437 (
    .I(seg_14_15_sp4_h_r_47_46977),
    .O(seg_14_15_local_g2_7_58396)
  );
  Span4Mux_h4 t1438 (
    .I(seg_11_15_sp4_v_t_40_43283),
    .O(seg_14_15_sp4_h_r_47_46977)
  );
  LocalMux t1439 (
    .I(seg_15_12_sp4_v_b_42_58116),
    .O(seg_15_12_local_g3_2_61860)
  );
  CascadeMux t144 (
    .I(net_42266),
    .O(net_42266_cascademuxed)
  );
  Span4Mux_v4 t1440 (
    .I(seg_15_15_sp4_h_l_42_46984),
    .O(seg_15_12_sp4_v_b_42_58116)
  );
  Span4Mux_h4 t1441 (
    .I(seg_11_15_sp4_v_t_42_43285),
    .O(seg_15_15_sp4_h_l_42_46984)
  );
  LocalMux t1442 (
    .I(seg_15_15_sp4_h_r_7_62306),
    .O(seg_15_15_local_g0_7_62210)
  );
  Span4Mux_h4 t1443 (
    .I(seg_15_15_sp4_h_l_42_46984),
    .O(seg_15_15_sp4_h_r_7_62306)
  );
  LocalMux t1444 (
    .I(seg_12_12_sp4_h_r_12_46607),
    .O(seg_12_12_local_g0_4_50347)
  );
  Span4Mux_h4 t1445 (
    .I(seg_11_12_sp4_v_t_45_42919),
    .O(seg_12_12_sp4_h_r_12_46607)
  );
  Span4Mux_v4 t1446 (
    .I(seg_11_16_sp4_v_t_37_43403),
    .O(seg_11_12_sp4_v_t_45_42919)
  );
  LocalMux t1447 (
    .I(seg_13_16_sp4_h_r_24_47098),
    .O(seg_13_16_local_g3_0_54690)
  );
  Span4Mux_h4 t1448 (
    .I(seg_11_16_sp4_v_t_37_43403),
    .O(seg_13_16_sp4_h_r_24_47098)
  );
  LocalMux t1449 (
    .I(seg_12_12_sp4_h_r_14_46611),
    .O(seg_12_12_local_g0_6_50349)
  );
  CascadeMux t145 (
    .I(net_42482),
    .O(net_42482_cascademuxed)
  );
  Span4Mux_h4 t1450 (
    .I(seg_11_12_sp4_v_t_47_42921),
    .O(seg_12_12_sp4_h_r_14_46611)
  );
  Span4Mux_v4 t1451 (
    .I(seg_11_16_sp4_v_t_39_43405),
    .O(seg_11_12_sp4_v_t_47_42921)
  );
  LocalMux t1452 (
    .I(seg_13_16_sp4_h_r_31_47107),
    .O(seg_13_16_local_g3_7_54697)
  );
  Span4Mux_h4 t1453 (
    .I(seg_11_16_sp4_v_t_39_43405),
    .O(seg_13_16_sp4_h_r_31_47107)
  );
  LocalMux t1454 (
    .I(seg_15_11_sp4_v_b_20_57749),
    .O(seg_15_11_local_g0_4_61715)
  );
  Span4Mux_v4 t1455 (
    .I(seg_15_12_sp4_h_l_38_46611),
    .O(seg_15_11_sp4_v_b_20_57749)
  );
  Span4Mux_h4 t1456 (
    .I(seg_11_12_sp4_v_t_47_42921),
    .O(seg_15_12_sp4_h_l_38_46611)
  );
  LocalMux t1457 (
    .I(seg_12_12_sp4_h_r_20_46617),
    .O(seg_12_12_local_g1_4_50355)
  );
  Span4Mux_h4 t1458 (
    .I(seg_11_12_sp4_v_t_41_42915),
    .O(seg_12_12_sp4_h_r_20_46617)
  );
  Span4Mux_v4 t1459 (
    .I(seg_11_16_sp4_v_t_41_43407),
    .O(seg_11_12_sp4_v_t_41_42915)
  );
  CascadeMux t146 (
    .I(net_42593),
    .O(net_42593_cascademuxed)
  );
  LocalMux t1460 (
    .I(seg_14_16_sp4_h_r_41_47104),
    .O(seg_14_16_local_g2_1_58513)
  );
  Span4Mux_h4 t1461 (
    .I(seg_11_16_sp4_v_t_41_43407),
    .O(seg_14_16_sp4_h_r_41_47104)
  );
  LocalMux t1462 (
    .I(seg_11_12_sp4_v_b_21_42550),
    .O(seg_11_12_local_g1_5_46525)
  );
  Span4Mux_v4 t1463 (
    .I(seg_11_13_sp4_v_t_40_43037),
    .O(seg_11_12_sp4_v_b_21_42550)
  );
  LocalMux t1464 (
    .I(seg_15_11_sp4_v_b_34_57875),
    .O(seg_15_11_local_g3_2_61737)
  );
  Span4Mux_v4 t1465 (
    .I(seg_15_13_sp4_h_l_47_46731),
    .O(seg_15_11_sp4_v_b_34_57875)
  );
  Span4Mux_h4 t1466 (
    .I(seg_11_13_sp4_v_t_40_43037),
    .O(seg_15_13_sp4_h_l_47_46731)
  );
  LocalMux t1467 (
    .I(seg_11_15_sp4_v_b_33_43041),
    .O(seg_11_15_local_g2_1_46898)
  );
  LocalMux t1468 (
    .I(seg_15_11_sp4_v_b_33_57872),
    .O(seg_15_11_local_g2_1_61728)
  );
  Span4Mux_v4 t1469 (
    .I(seg_15_13_sp4_h_l_44_46740),
    .O(seg_15_11_sp4_v_b_33_57872)
  );
  CascadeMux t147 (
    .I(net_42605),
    .O(net_42605_cascademuxed)
  );
  Span4Mux_h4 t1470 (
    .I(seg_11_13_sp4_v_t_44_43041),
    .O(seg_15_13_sp4_h_l_44_46740)
  );
  LocalMux t1471 (
    .I(seg_10_12_sp4_v_b_23_38721),
    .O(seg_10_12_local_g1_7_42696)
  );
  Span4Mux_v4 t1472 (
    .I(seg_10_13_sp4_v_t_47_39213),
    .O(seg_10_12_sp4_v_b_23_38721)
  );
  LocalMux t1473 (
    .I(seg_10_12_sp4_v_b_25_38833),
    .O(seg_10_12_local_g2_1_42698)
  );
  Span4Mux_v4 t1474 (
    .I(seg_10_14_sp4_v_t_36_39325),
    .O(seg_10_12_sp4_v_b_25_38833)
  );
  LocalMux t1475 (
    .I(seg_10_14_sp4_h_r_8_43031),
    .O(seg_10_14_local_g0_0_42927)
  );
  Span4Mux_h4 t1476 (
    .I(seg_10_14_sp4_v_t_38_39327),
    .O(seg_10_14_sp4_h_r_8_43031)
  );
  LocalMux t1477 (
    .I(seg_10_13_sp4_v_b_26_38959),
    .O(seg_10_13_local_g2_2_42822)
  );
  Span4Mux_v4 t1478 (
    .I(seg_10_15_sp4_v_t_43_39455),
    .O(seg_10_13_sp4_v_b_26_38959)
  );
  LocalMux t1479 (
    .I(seg_10_12_sp4_v_b_13_38711),
    .O(seg_10_12_local_g0_5_42686)
  );
  CascadeMux t148 (
    .I(net_42716),
    .O(net_42716_cascademuxed)
  );
  Span4Mux_v4 t1480 (
    .I(seg_10_13_sp4_v_t_41_39207),
    .O(seg_10_12_sp4_v_b_13_38711)
  );
  LocalMux t1481 (
    .I(seg_13_12_sp4_r_v_b_23_54045),
    .O(seg_13_12_local_g3_7_54205)
  );
  Span4Mux_v4 t1482 (
    .I(seg_14_13_sp4_h_l_41_42904),
    .O(seg_13_12_sp4_r_v_b_23_54045)
  );
  Span4Mux_h4 t1483 (
    .I(seg_10_13_sp4_v_t_41_39207),
    .O(seg_14_13_sp4_h_l_41_42904)
  );
  LocalMux t1484 (
    .I(seg_13_16_sp4_h_r_37_43267),
    .O(seg_13_16_local_g2_5_54687)
  );
  Span4Mux_h4 t1485 (
    .I(seg_10_16_sp4_v_t_42_39577),
    .O(seg_13_16_sp4_h_r_37_43267)
  );
  LocalMux t1486 (
    .I(seg_13_16_sp4_h_r_44_43278),
    .O(seg_13_16_local_g3_4_54694)
  );
  Span4Mux_h4 t1487 (
    .I(seg_10_16_sp4_v_t_44_39579),
    .O(seg_13_16_sp4_h_r_44_43278)
  );
  LocalMux t1488 (
    .I(seg_10_12_sp4_v_b_20_38718),
    .O(seg_10_12_local_g0_4_42685)
  );
  Span4Mux_v4 t1489 (
    .I(seg_10_13_sp4_v_t_43_39209),
    .O(seg_10_12_sp4_v_b_20_38718)
  );
  CascadeMux t149 (
    .I(net_42722),
    .O(net_42722_cascademuxed)
  );
  LocalMux t1490 (
    .I(seg_13_13_sp4_h_r_46_42901),
    .O(seg_13_13_local_g2_6_54319)
  );
  Span4Mux_h4 t1491 (
    .I(seg_10_13_sp4_v_t_43_39209),
    .O(seg_13_13_sp4_h_r_46_42901)
  );
  LocalMux t1492 (
    .I(seg_10_12_sp4_v_b_22_38720),
    .O(seg_10_12_local_g0_6_42687)
  );
  Span4Mux_v4 t1493 (
    .I(seg_10_13_sp4_v_t_45_39211),
    .O(seg_10_12_sp4_v_b_22_38720)
  );
  LocalMux t1494 (
    .I(seg_10_15_sp4_v_b_32_39211),
    .O(seg_10_15_local_g3_0_43074)
  );
  LocalMux t1495 (
    .I(seg_10_18_lutff_0_out_39547),
    .O(seg_10_18_local_g3_0_43443)
  );
  LocalMux t1496 (
    .I(seg_10_18_lutff_1_out_39548),
    .O(seg_10_18_local_g2_1_43436)
  );
  LocalMux t1497 (
    .I(seg_10_18_lutff_2_out_39549),
    .O(seg_10_18_local_g2_2_43437)
  );
  LocalMux t1498 (
    .I(seg_10_18_lutff_3_out_39550),
    .O(seg_10_18_local_g1_3_43430)
  );
  LocalMux t1499 (
    .I(seg_10_18_lutff_4_out_39551),
    .O(seg_10_18_local_g3_4_43447)
  );
  CascadeMux t15 (
    .I(net_13560),
    .O(net_13560_cascademuxed)
  );
  CascadeMux t150 (
    .I(net_42728),
    .O(net_42728_cascademuxed)
  );
  LocalMux t1500 (
    .I(seg_10_18_lutff_5_out_39552),
    .O(seg_10_18_local_g0_5_43424)
  );
  LocalMux t1501 (
    .I(seg_10_18_lutff_6_out_39553),
    .O(seg_10_18_local_g2_6_43441)
  );
  LocalMux t1502 (
    .I(seg_10_18_lutff_7_out_39554),
    .O(seg_10_18_local_g3_7_43450)
  );
  LocalMux t1503 (
    .I(seg_15_18_sp4_h_r_35_55009),
    .O(seg_15_18_local_g3_3_62599)
  );
  Span4Mux_h4 t1504 (
    .I(seg_13_18_sp4_h_l_38_39687),
    .O(seg_15_18_sp4_h_r_35_55009)
  );
  LocalMux t1505 (
    .I(seg_16_18_sp4_h_r_46_55009),
    .O(seg_16_18_local_g3_6_66433)
  );
  Span4Mux_h4 t1506 (
    .I(seg_13_18_sp4_h_l_38_39687),
    .O(seg_16_18_sp4_h_r_46_55009)
  );
  LocalMux t1507 (
    .I(seg_12_13_sp4_r_v_b_21_50335),
    .O(seg_12_13_local_g3_5_50495)
  );
  Span4Mux_v4 t1508 (
    .I(seg_13_14_sp4_v_t_40_50822),
    .O(seg_12_13_sp4_r_v_b_21_50335)
  );
  Span4Mux_v4 t1509 (
    .I(seg_13_18_sp4_h_l_40_39689),
    .O(seg_13_14_sp4_v_t_40_50822)
  );
  CascadeMux t151 (
    .I(net_42734),
    .O(net_42734_cascademuxed)
  );
  LocalMux t1510 (
    .I(seg_13_17_sp4_v_b_16_50822),
    .O(seg_13_17_local_g0_0_54789)
  );
  Span4Mux_v4 t1511 (
    .I(seg_13_18_sp4_h_l_40_39689),
    .O(seg_13_17_sp4_v_b_16_50822)
  );
  LocalMux t1512 (
    .I(seg_13_17_sp4_v_b_12_50818),
    .O(seg_13_17_local_g1_4_54801)
  );
  Span4Mux_v4 t1513 (
    .I(seg_13_18_sp4_h_l_42_39691),
    .O(seg_13_17_sp4_v_b_12_50818)
  );
  LocalMux t1514 (
    .I(seg_12_16_sp4_r_v_b_35_50828),
    .O(seg_12_16_local_g2_3_50854)
  );
  Span4Mux_v4 t1515 (
    .I(seg_13_18_sp4_h_l_46_39685),
    .O(seg_12_16_sp4_r_v_b_35_50828)
  );
  LocalMux t1516 (
    .I(seg_12_13_sp4_v_b_15_46498),
    .O(seg_12_13_local_g1_7_50481)
  );
  Span4Mux_v4 t1517 (
    .I(seg_12_14_sp4_v_t_43_46994),
    .O(seg_12_13_sp4_v_b_15_46498)
  );
  Span4Mux_v4 t1518 (
    .I(seg_12_18_sp4_h_l_37_35851),
    .O(seg_12_14_sp4_v_t_43_46994)
  );
  LocalMux t1519 (
    .I(seg_12_16_sp4_v_b_30_46994),
    .O(seg_12_16_local_g3_6_50865)
  );
  CascadeMux t152 (
    .I(net_42740),
    .O(net_42740_cascademuxed)
  );
  Span4Mux_v4 t1520 (
    .I(seg_12_18_sp4_h_l_37_35851),
    .O(seg_12_16_sp4_v_b_30_46994)
  );
  LocalMux t1521 (
    .I(seg_12_13_sp4_v_b_17_46500),
    .O(seg_12_13_local_g0_1_50467)
  );
  Span4Mux_v4 t1522 (
    .I(seg_12_14_sp4_v_t_45_46996),
    .O(seg_12_13_sp4_v_b_17_46500)
  );
  Span4Mux_v4 t1523 (
    .I(seg_12_18_sp4_h_l_39_35855),
    .O(seg_12_14_sp4_v_t_45_46996)
  );
  LocalMux t1524 (
    .I(seg_15_17_sp4_r_v_b_22_62319),
    .O(seg_15_17_local_g3_6_62479)
  );
  Span4Mux_v4 t1525 (
    .I(seg_16_18_sp4_h_l_46_51178),
    .O(seg_15_17_sp4_r_v_b_22_62319)
  );
  Span4Mux_h4 t1526 (
    .I(seg_12_18_sp4_h_l_45_35861),
    .O(seg_16_18_sp4_h_l_46_51178)
  );
  LocalMux t1527 (
    .I(seg_12_13_sp4_v_b_12_46495),
    .O(seg_12_13_local_g1_4_50478)
  );
  Span4Mux_v4 t1528 (
    .I(seg_12_14_sp4_v_t_47_46998),
    .O(seg_12_13_sp4_v_b_12_46495)
  );
  Span4Mux_v4 t1529 (
    .I(seg_12_18_sp4_h_l_47_35853),
    .O(seg_12_14_sp4_v_t_47_46998)
  );
  CascadeMux t153 (
    .I(net_42746),
    .O(net_42746_cascademuxed)
  );
  LocalMux t1530 (
    .I(seg_15_17_sp4_r_v_b_12_62309),
    .O(seg_15_17_local_g2_4_62469)
  );
  Span4Mux_v4 t1531 (
    .I(seg_16_18_sp4_h_l_36_51176),
    .O(seg_15_17_sp4_r_v_b_12_62309)
  );
  Span4Mux_h4 t1532 (
    .I(seg_12_18_sp4_h_l_47_35853),
    .O(seg_16_18_sp4_h_l_36_51176)
  );
  LocalMux t1533 (
    .I(seg_13_17_sp4_r_v_b_17_54654),
    .O(seg_13_17_local_g3_1_54814)
  );
  Span4Mux_v4 t1534 (
    .I(seg_14_18_sp4_h_l_41_43519),
    .O(seg_13_17_sp4_r_v_b_17_54654)
  );
  LocalMux t1535 (
    .I(seg_14_17_sp4_v_b_17_54654),
    .O(seg_14_17_local_g0_1_58620)
  );
  Span4Mux_v4 t1536 (
    .I(seg_14_18_sp4_h_l_41_43519),
    .O(seg_14_17_sp4_v_b_17_54654)
  );
  LocalMux t1537 (
    .I(seg_13_17_sp4_r_v_b_21_54658),
    .O(seg_13_17_local_g3_5_54818)
  );
  Span4Mux_v4 t1538 (
    .I(seg_14_18_sp4_h_l_45_43523),
    .O(seg_13_17_sp4_r_v_b_21_54658)
  );
  LocalMux t1539 (
    .I(seg_11_12_sp4_v_b_28_42669),
    .O(seg_11_12_local_g2_4_46532)
  );
  CascadeMux t154 (
    .I(net_42752),
    .O(net_42752_cascademuxed)
  );
  Span4Mux_v4 t1540 (
    .I(seg_11_14_sp4_v_t_36_43156),
    .O(seg_11_12_sp4_v_b_28_42669)
  );
  LocalMux t1541 (
    .I(seg_14_13_sp4_r_v_b_12_57987),
    .O(seg_14_13_local_g2_4_58147)
  );
  Span4Mux_v4 t1542 (
    .I(seg_15_14_sp4_h_l_36_46853),
    .O(seg_14_13_sp4_r_v_b_12_57987)
  );
  Span4Mux_h4 t1543 (
    .I(seg_11_14_sp4_v_t_36_43156),
    .O(seg_15_14_sp4_h_l_36_46853)
  );
  LocalMux t1544 (
    .I(seg_15_12_sp4_v_b_25_57987),
    .O(seg_15_12_local_g2_1_61851)
  );
  Span4Mux_v4 t1545 (
    .I(seg_15_14_sp4_h_l_36_46853),
    .O(seg_15_12_sp4_v_b_25_57987)
  );
  LocalMux t1546 (
    .I(seg_15_14_sp4_v_b_1_57987),
    .O(seg_15_14_local_g0_1_62081)
  );
  Span4Mux_v4 t1547 (
    .I(seg_15_14_sp4_h_l_36_46853),
    .O(seg_15_14_sp4_v_b_1_57987)
  );
  LocalMux t1548 (
    .I(seg_13_14_sp4_h_r_35_46855),
    .O(seg_13_14_local_g3_3_54447)
  );
  Span4Mux_h4 t1549 (
    .I(seg_11_14_sp4_v_t_46_43166),
    .O(seg_13_14_sp4_h_r_35_46855)
  );
  CascadeMux t155 (
    .I(net_42758),
    .O(net_42758_cascademuxed)
  );
  LocalMux t1550 (
    .I(seg_15_12_sp4_v_b_29_57991),
    .O(seg_15_12_local_g3_5_61863)
  );
  Span4Mux_v4 t1551 (
    .I(seg_15_14_sp4_h_l_46_46855),
    .O(seg_15_12_sp4_v_b_29_57991)
  );
  Span4Mux_h4 t1552 (
    .I(seg_11_14_sp4_v_t_46_43166),
    .O(seg_15_14_sp4_h_l_46_46855)
  );
  LocalMux t1553 (
    .I(seg_11_15_sp4_h_r_5_46982),
    .O(seg_11_15_local_g1_5_46894)
  );
  Span4Mux_h4 t1554 (
    .I(seg_11_15_sp4_v_t_37_43280),
    .O(seg_11_15_sp4_h_r_5_46982)
  );
  LocalMux t1555 (
    .I(seg_12_15_sp4_h_r_16_46982),
    .O(seg_12_15_local_g0_0_50712)
  );
  Span4Mux_h4 t1556 (
    .I(seg_11_15_sp4_v_t_37_43280),
    .O(seg_12_15_sp4_h_r_16_46982)
  );
  LocalMux t1557 (
    .I(seg_13_15_sp4_h_r_29_46982),
    .O(seg_13_15_local_g2_5_54564)
  );
  Span4Mux_h4 t1558 (
    .I(seg_11_15_sp4_v_t_37_43280),
    .O(seg_13_15_sp4_h_r_29_46982)
  );
  LocalMux t1559 (
    .I(seg_15_12_sp4_v_b_46_58120),
    .O(seg_15_12_local_g3_6_61864)
  );
  CascadeMux t156 (
    .I(net_42839),
    .O(net_42839_cascademuxed)
  );
  Span4Mux_v4 t1560 (
    .I(seg_15_15_sp4_h_l_40_46982),
    .O(seg_15_12_sp4_v_b_46_58120)
  );
  Span4Mux_h4 t1561 (
    .I(seg_11_15_sp4_v_t_37_43280),
    .O(seg_15_15_sp4_h_l_40_46982)
  );
  LocalMux t1562 (
    .I(seg_16_19_sp4_h_r_17_62795),
    .O(seg_16_19_local_g0_1_66527)
  );
  Span4Mux_h4 t1563 (
    .I(seg_15_19_sp4_h_l_45_47477),
    .O(seg_16_19_sp4_h_r_17_62795)
  );
  Span4Mux_h4 t1564 (
    .I(seg_11_19_sp4_v_b_2_43282),
    .O(seg_15_19_sp4_h_l_45_47477)
  );
  LocalMux t1565 (
    .I(seg_15_12_sp4_v_b_40_58114),
    .O(seg_15_12_local_g2_0_61850)
  );
  Span4Mux_v4 t1566 (
    .I(seg_15_15_sp4_h_l_46_46978),
    .O(seg_15_12_sp4_v_b_40_58114)
  );
  Span4Mux_h4 t1567 (
    .I(seg_11_15_sp4_v_t_43_43286),
    .O(seg_15_15_sp4_h_l_46_46978)
  );
  LocalMux t1568 (
    .I(seg_11_15_sp4_h_r_3_46980),
    .O(seg_11_15_local_g0_3_46884)
  );
  Span4Mux_h4 t1569 (
    .I(seg_11_15_sp4_v_t_47_43290),
    .O(seg_11_15_sp4_h_r_3_46980)
  );
  CascadeMux t157 (
    .I(net_42845),
    .O(net_42845_cascademuxed)
  );
  LocalMux t1570 (
    .I(seg_12_15_sp4_h_r_14_46980),
    .O(seg_12_15_local_g1_6_50726)
  );
  Span4Mux_h4 t1571 (
    .I(seg_11_15_sp4_v_t_47_43290),
    .O(seg_12_15_sp4_h_r_14_46980)
  );
  LocalMux t1572 (
    .I(seg_13_15_sp4_h_r_27_46980),
    .O(seg_13_15_local_g2_3_54562)
  );
  Span4Mux_h4 t1573 (
    .I(seg_11_15_sp4_v_t_47_43290),
    .O(seg_13_15_sp4_h_r_27_46980)
  );
  LocalMux t1574 (
    .I(seg_15_12_sp4_v_b_38_58112),
    .O(seg_15_12_local_g2_6_61856)
  );
  Span4Mux_v4 t1575 (
    .I(seg_15_15_sp4_h_l_38_46980),
    .O(seg_15_12_sp4_v_b_38_58112)
  );
  Span4Mux_h4 t1576 (
    .I(seg_11_15_sp4_v_t_47_43290),
    .O(seg_15_15_sp4_h_l_38_46980)
  );
  LocalMux t1577 (
    .I(seg_11_14_sp4_h_r_8_46862),
    .O(seg_11_14_local_g0_0_46758)
  );
  Span4Mux_h4 t1578 (
    .I(seg_11_14_sp4_v_t_38_43158),
    .O(seg_11_14_sp4_h_r_8_46862)
  );
  LocalMux t1579 (
    .I(seg_15_14_sp4_h_r_11_62177),
    .O(seg_15_14_local_g0_3_62083)
  );
  CascadeMux t158 (
    .I(net_42851),
    .O(net_42851_cascademuxed)
  );
  Span4Mux_h4 t1580 (
    .I(seg_15_14_sp4_h_l_45_46862),
    .O(seg_15_14_sp4_h_r_11_62177)
  );
  Span4Mux_h4 t1581 (
    .I(seg_11_14_sp4_v_t_38_43158),
    .O(seg_15_14_sp4_h_l_45_46862)
  );
  LocalMux t1582 (
    .I(seg_16_20_sp4_h_r_20_62923),
    .O(seg_16_20_local_g1_4_66661)
  );
  Span4Mux_h4 t1583 (
    .I(seg_15_20_sp4_h_l_36_47591),
    .O(seg_16_20_sp4_h_r_20_62923)
  );
  Span4Mux_h4 t1584 (
    .I(seg_11_20_sp4_v_b_7_43408),
    .O(seg_15_20_sp4_h_l_36_47591)
  );
  LocalMux t1585 (
    .I(seg_12_13_sp4_h_r_16_46736),
    .O(seg_12_13_local_g0_0_50466)
  );
  Span4Mux_h4 t1586 (
    .I(seg_11_13_sp4_v_t_37_43034),
    .O(seg_12_13_sp4_h_r_16_46736)
  );
  Span4Mux_v4 t1587 (
    .I(seg_11_17_sp4_v_t_37_43526),
    .O(seg_11_13_sp4_v_t_37_43034)
  );
  LocalMux t1588 (
    .I(seg_12_13_sp4_h_r_18_46738),
    .O(seg_12_13_local_g0_2_50468)
  );
  Span4Mux_h4 t1589 (
    .I(seg_11_13_sp4_v_t_39_43036),
    .O(seg_12_13_sp4_h_r_18_46738)
  );
  CascadeMux t159 (
    .I(net_42857),
    .O(net_42857_cascademuxed)
  );
  Span4Mux_v4 t1590 (
    .I(seg_11_17_sp4_v_t_39_43528),
    .O(seg_11_13_sp4_v_t_39_43036)
  );
  LocalMux t1591 (
    .I(seg_13_17_sp4_h_r_31_47230),
    .O(seg_13_17_local_g3_7_54820)
  );
  Span4Mux_h4 t1592 (
    .I(seg_11_17_sp4_v_t_39_43528),
    .O(seg_13_17_sp4_h_r_31_47230)
  );
  LocalMux t1593 (
    .I(seg_13_17_sp4_h_r_30_47229),
    .O(seg_13_17_local_g2_6_54811)
  );
  Span4Mux_h4 t1594 (
    .I(seg_11_17_sp4_v_t_43_43532),
    .O(seg_13_17_sp4_h_r_30_47229)
  );
  LocalMux t1595 (
    .I(seg_15_15_sp4_v_b_35_58366),
    .O(seg_15_15_local_g3_3_62230)
  );
  Span4Mux_v4 t1596 (
    .I(seg_15_17_sp4_h_l_46_47224),
    .O(seg_15_15_sp4_v_b_35_58366)
  );
  Span4Mux_h4 t1597 (
    .I(seg_11_17_sp4_v_t_43_43532),
    .O(seg_15_17_sp4_h_l_46_47224)
  );
  LocalMux t1598 (
    .I(seg_15_17_sp4_h_r_7_62552),
    .O(seg_15_17_local_g0_7_62456)
  );
  Span4Mux_h4 t1599 (
    .I(seg_15_17_sp4_h_l_46_47224),
    .O(seg_15_17_sp4_h_r_7_62552)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t16 (
    .carryinitin(net_17430),
    .carryinitout(net_17474)
  );
  CascadeMux t160 (
    .I(net_42863),
    .O(net_42863_cascademuxed)
  );
  LocalMux t1600 (
    .I(seg_12_13_sp4_h_r_21_46739),
    .O(seg_12_13_local_g0_5_50471)
  );
  Span4Mux_h4 t1601 (
    .I(seg_11_13_sp4_v_t_45_43042),
    .O(seg_12_13_sp4_h_r_21_46739)
  );
  Span4Mux_v4 t1602 (
    .I(seg_11_17_sp4_v_t_45_43534),
    .O(seg_11_13_sp4_v_t_45_43042)
  );
  LocalMux t1603 (
    .I(seg_12_17_sp4_h_r_21_47231),
    .O(seg_12_17_local_g0_5_50963)
  );
  Span4Mux_h4 t1604 (
    .I(seg_11_17_sp4_v_t_45_43534),
    .O(seg_12_17_sp4_h_r_21_47231)
  );
  LocalMux t1605 (
    .I(seg_13_17_sp4_h_r_32_47231),
    .O(seg_13_17_local_g2_0_54805)
  );
  Span4Mux_h4 t1606 (
    .I(seg_11_17_sp4_v_t_45_43534),
    .O(seg_13_17_sp4_h_r_32_47231)
  );
  LocalMux t1607 (
    .I(seg_11_14_sp4_h_r_10_46854),
    .O(seg_11_14_local_g0_2_46760)
  );
  Span4Mux_h4 t1608 (
    .I(seg_11_14_sp4_v_t_40_43160),
    .O(seg_11_14_sp4_h_r_10_46854)
  );
  LocalMux t1609 (
    .I(seg_14_14_sp4_h_r_40_46859),
    .O(seg_14_14_local_g3_0_58274)
  );
  CascadeMux t161 (
    .I(net_42869),
    .O(net_42869_cascademuxed)
  );
  Span4Mux_h4 t1610 (
    .I(seg_11_14_sp4_v_t_40_43160),
    .O(seg_14_14_sp4_h_r_40_46859)
  );
  LocalMux t1611 (
    .I(seg_15_12_sp4_v_b_34_57998),
    .O(seg_15_12_local_g2_2_61852)
  );
  Span4Mux_v4 t1612 (
    .I(seg_15_14_sp4_h_l_47_46854),
    .O(seg_15_12_sp4_v_b_34_57998)
  );
  Span4Mux_h4 t1613 (
    .I(seg_11_14_sp4_v_t_40_43160),
    .O(seg_15_14_sp4_h_l_47_46854)
  );
  LocalMux t1614 (
    .I(seg_13_14_sp4_h_r_33_46863),
    .O(seg_13_14_local_g2_1_54437)
  );
  Span4Mux_h4 t1615 (
    .I(seg_11_14_sp4_v_t_44_43164),
    .O(seg_13_14_sp4_h_r_33_46863)
  );
  LocalMux t1616 (
    .I(seg_14_14_sp4_h_r_44_46863),
    .O(seg_14_14_local_g2_4_58270)
  );
  Span4Mux_h4 t1617 (
    .I(seg_11_14_sp4_v_t_44_43164),
    .O(seg_14_14_sp4_h_r_44_46863)
  );
  LocalMux t1618 (
    .I(seg_15_12_sp4_v_b_27_57989),
    .O(seg_15_12_local_g3_3_61861)
  );
  Span4Mux_v4 t1619 (
    .I(seg_15_14_sp4_h_l_44_46863),
    .O(seg_15_12_sp4_v_b_27_57989)
  );
  CascadeMux t162 (
    .I(net_42875),
    .O(net_42875_cascademuxed)
  );
  Span4Mux_h4 t1620 (
    .I(seg_11_14_sp4_v_t_44_43164),
    .O(seg_15_14_sp4_h_l_44_46863)
  );
  LocalMux t1621 (
    .I(seg_10_13_sp4_v_b_21_38842),
    .O(seg_10_13_local_g0_5_42809)
  );
  Span4Mux_v4 t1622 (
    .I(seg_10_14_sp4_v_t_37_39326),
    .O(seg_10_13_sp4_v_b_21_38842)
  );
  LocalMux t1623 (
    .I(seg_10_13_sp4_v_b_19_38840),
    .O(seg_10_13_local_g1_3_42815)
  );
  Span4Mux_v4 t1624 (
    .I(seg_10_14_sp4_v_t_47_39336),
    .O(seg_10_13_sp4_v_b_19_38840)
  );
  LocalMux t1625 (
    .I(seg_13_13_sp4_r_v_b_23_54168),
    .O(seg_13_13_local_g3_7_54328)
  );
  Span4Mux_v4 t1626 (
    .I(seg_14_14_sp4_h_l_47_43023),
    .O(seg_13_13_sp4_r_v_b_23_54168)
  );
  Span4Mux_h4 t1627 (
    .I(seg_10_14_sp4_v_t_47_39336),
    .O(seg_14_14_sp4_h_l_47_43023)
  );
  LocalMux t1628 (
    .I(seg_10_13_sp4_v_b_28_38961),
    .O(seg_10_13_local_g3_4_42832)
  );
  Span4Mux_v4 t1629 (
    .I(seg_10_15_sp4_v_t_36_39448),
    .O(seg_10_13_sp4_v_b_28_38961)
  );
  CascadeMux t163 (
    .I(net_42881),
    .O(net_42881_cascademuxed)
  );
  LocalMux t1630 (
    .I(seg_10_13_sp4_v_b_16_38837),
    .O(seg_10_13_local_g0_0_42804)
  );
  Span4Mux_v4 t1631 (
    .I(seg_10_14_sp4_v_t_39_39328),
    .O(seg_10_13_sp4_v_b_16_38837)
  );
  LocalMux t1632 (
    .I(seg_10_14_sp4_h_r_7_43030),
    .O(seg_10_14_local_g1_7_42942)
  );
  Span4Mux_h4 t1633 (
    .I(seg_10_14_sp4_v_t_39_39328),
    .O(seg_10_14_sp4_h_r_7_43030)
  );
  LocalMux t1634 (
    .I(seg_10_13_sp4_v_b_13_38834),
    .O(seg_10_13_local_g1_5_42817)
  );
  Span4Mux_v4 t1635 (
    .I(seg_10_14_sp4_v_t_41_39330),
    .O(seg_10_13_sp4_v_b_13_38834)
  );
  LocalMux t1636 (
    .I(seg_10_14_sp4_h_r_9_43032),
    .O(seg_10_14_local_g1_1_42936)
  );
  Span4Mux_h4 t1637 (
    .I(seg_10_14_sp4_v_t_41_39330),
    .O(seg_10_14_sp4_h_r_9_43032)
  );
  LocalMux t1638 (
    .I(seg_10_13_sp4_v_b_20_38841),
    .O(seg_10_13_local_g0_4_42808)
  );
  Span4Mux_v4 t1639 (
    .I(seg_10_14_sp4_v_t_43_39332),
    .O(seg_10_13_sp4_v_b_20_38841)
  );
  CascadeMux t164 (
    .I(net_42962),
    .O(net_42962_cascademuxed)
  );
  LocalMux t1640 (
    .I(seg_10_13_sp4_v_b_17_38838),
    .O(seg_10_13_local_g1_1_42813)
  );
  Span4Mux_v4 t1641 (
    .I(seg_10_14_sp4_v_t_45_39334),
    .O(seg_10_13_sp4_v_b_17_38838)
  );
  LocalMux t1642 (
    .I(seg_13_13_sp4_r_v_b_18_54163),
    .O(seg_13_13_local_g3_2_54323)
  );
  Span4Mux_v4 t1643 (
    .I(seg_14_14_sp4_h_l_36_43022),
    .O(seg_13_13_sp4_r_v_b_18_54163)
  );
  Span4Mux_h4 t1644 (
    .I(seg_10_14_sp4_v_t_45_39334),
    .O(seg_14_14_sp4_h_l_36_43022)
  );
  LocalMux t1645 (
    .I(seg_10_19_lutff_0_out_39670),
    .O(seg_10_19_local_g1_0_43550)
  );
  LocalMux t1646 (
    .I(seg_11_18_neigh_op_tnl_0_39670),
    .O(seg_11_18_local_g3_0_47274)
  );
  LocalMux t1647 (
    .I(seg_10_19_lutff_1_out_39671),
    .O(seg_10_19_local_g1_1_43551)
  );
  LocalMux t1648 (
    .I(seg_11_19_neigh_op_lft_1_39671),
    .O(seg_11_19_local_g0_1_47374)
  );
  LocalMux t1649 (
    .I(seg_10_19_lutff_2_out_39672),
    .O(seg_10_19_local_g0_2_43544)
  );
  CascadeMux t165 (
    .I(net_42974),
    .O(net_42974_cascademuxed)
  );
  LocalMux t1650 (
    .I(seg_10_19_lutff_3_out_39673),
    .O(seg_10_19_local_g3_3_43569)
  );
  LocalMux t1651 (
    .I(seg_10_19_lutff_4_out_39674),
    .O(seg_10_19_local_g1_4_43554)
  );
  LocalMux t1652 (
    .I(seg_11_19_neigh_op_lft_4_39674),
    .O(seg_11_19_local_g1_4_47385)
  );
  LocalMux t1653 (
    .I(seg_11_20_neigh_op_bnl_4_39674),
    .O(seg_11_20_local_g2_4_47516)
  );
  LocalMux t1654 (
    .I(seg_9_18_neigh_op_tnr_5_39675),
    .O(seg_9_18_local_g2_5_39609)
  );
  LocalMux t1655 (
    .I(seg_10_19_lutff_5_out_39675),
    .O(seg_10_19_local_g3_5_43571)
  );
  LocalMux t1656 (
    .I(seg_11_18_neigh_op_tnl_5_39675),
    .O(seg_11_18_local_g3_5_47279)
  );
  LocalMux t1657 (
    .I(seg_9_18_neigh_op_tnr_6_39676),
    .O(seg_9_18_local_g2_6_39610)
  );
  LocalMux t1658 (
    .I(seg_10_19_lutff_6_out_39676),
    .O(seg_10_19_local_g0_6_43548)
  );
  LocalMux t1659 (
    .I(seg_11_18_neigh_op_tnl_6_39676),
    .O(seg_11_18_local_g2_6_47272)
  );
  CascadeMux t166 (
    .I(net_42992),
    .O(net_42992_cascademuxed)
  );
  LocalMux t1660 (
    .I(seg_10_19_lutff_7_out_39677),
    .O(seg_10_19_local_g0_7_43549)
  );
  LocalMux t1661 (
    .I(seg_12_19_sp4_h_r_24_43636),
    .O(seg_12_19_local_g2_0_51220)
  );
  LocalMux t1662 (
    .I(seg_13_18_sp4_r_v_b_13_54773),
    .O(seg_13_18_local_g2_5_54933)
  );
  Span4Mux_v4 t1663 (
    .I(seg_14_19_sp4_h_l_37_43636),
    .O(seg_13_18_sp4_r_v_b_13_54773)
  );
  LocalMux t1664 (
    .I(seg_13_18_sp4_r_v_b_23_54783),
    .O(seg_13_18_local_g3_7_54943)
  );
  Span4Mux_v4 t1665 (
    .I(seg_14_19_sp4_h_l_47_43638),
    .O(seg_13_18_sp4_r_v_b_23_54783)
  );
  LocalMux t1666 (
    .I(seg_14_18_sp4_v_b_23_54783),
    .O(seg_14_18_local_g0_7_58749)
  );
  Span4Mux_v4 t1667 (
    .I(seg_14_19_sp4_h_l_47_43638),
    .O(seg_14_18_sp4_v_b_23_54783)
  );
  LocalMux t1668 (
    .I(seg_15_19_sp4_h_r_28_55135),
    .O(seg_15_19_local_g2_4_62715)
  );
  Span4Mux_h4 t1669 (
    .I(seg_13_19_sp4_h_l_36_39806),
    .O(seg_15_19_sp4_h_r_28_55135)
  );
  CascadeMux t167 (
    .I(net_42998),
    .O(net_42998_cascademuxed)
  );
  LocalMux t1670 (
    .I(seg_16_19_sp4_h_r_43_55137),
    .O(seg_16_19_local_g3_3_66553)
  );
  Span4Mux_h4 t1671 (
    .I(seg_13_19_sp4_h_l_38_39810),
    .O(seg_16_19_sp4_h_r_43_55137)
  );
  LocalMux t1672 (
    .I(seg_16_20_sp4_r_v_b_43_66762),
    .O(seg_16_20_local_g3_3_66676)
  );
  Span4Mux_v4 t1673 (
    .I(seg_17_19_sp4_h_l_43_55137),
    .O(seg_16_20_sp4_r_v_b_43_66762)
  );
  Span4Mux_h4 t1674 (
    .I(seg_13_19_sp4_h_l_38_39810),
    .O(seg_17_19_sp4_h_l_43_55137)
  );
  LocalMux t1675 (
    .I(seg_17_19_sp4_h_r_6_70459),
    .O(seg_17_19_local_g1_6_70371)
  );
  Span4Mux_h4 t1676 (
    .I(seg_17_19_sp4_h_l_43_55137),
    .O(seg_17_19_sp4_h_r_6_70459)
  );
  LocalMux t1677 (
    .I(seg_17_20_sp4_v_b_43_66762),
    .O(seg_17_20_local_g3_3_70507)
  );
  Span4Mux_v4 t1678 (
    .I(seg_17_19_sp4_h_l_43_55137),
    .O(seg_17_20_sp4_v_b_43_66762)
  );
  LocalMux t1679 (
    .I(seg_12_18_sp4_r_v_b_16_50945),
    .O(seg_12_18_local_g3_0_51105)
  );
  CascadeMux t168 (
    .I(net_43085),
    .O(net_43085_cascademuxed)
  );
  Span4Mux_v4 t1680 (
    .I(seg_13_19_sp4_h_l_40_39812),
    .O(seg_12_18_sp4_r_v_b_16_50945)
  );
  LocalMux t1681 (
    .I(seg_14_19_sp4_h_r_10_58961),
    .O(seg_14_19_local_g1_2_58875)
  );
  Span4Mux_h4 t1682 (
    .I(seg_14_19_sp4_h_l_39_43640),
    .O(seg_14_19_sp4_h_r_10_58961)
  );
  LocalMux t1683 (
    .I(seg_15_19_sp4_h_r_23_58961),
    .O(seg_15_19_local_g0_7_62702)
  );
  Span4Mux_h4 t1684 (
    .I(seg_14_19_sp4_h_l_39_43640),
    .O(seg_15_19_sp4_h_r_23_58961)
  );
  LocalMux t1685 (
    .I(seg_12_18_sp4_r_v_b_14_50943),
    .O(seg_12_18_local_g2_6_51103)
  );
  Span4Mux_v4 t1686 (
    .I(seg_13_19_sp4_h_l_44_39816),
    .O(seg_12_18_sp4_r_v_b_14_50943)
  );
  LocalMux t1687 (
    .I(seg_12_20_sp4_v_b_40_47606),
    .O(seg_12_20_local_g2_0_51343)
  );
  Span4Mux_v4 t1688 (
    .I(seg_12_19_sp4_h_l_37_35974),
    .O(seg_12_20_sp4_v_b_40_47606)
  );
  LocalMux t1689 (
    .I(seg_15_18_sp4_r_v_b_13_62433),
    .O(seg_15_18_local_g2_5_62593)
  );
  CascadeMux t169 (
    .I(net_43109),
    .O(net_43109_cascademuxed)
  );
  Span4Mux_v4 t1690 (
    .I(seg_16_19_sp4_h_l_37_51298),
    .O(seg_15_18_sp4_r_v_b_13_62433)
  );
  Span4Mux_h4 t1691 (
    .I(seg_12_19_sp4_h_l_41_35980),
    .O(seg_16_19_sp4_h_l_37_51298)
  );
  LocalMux t1692 (
    .I(seg_15_18_sp4_r_v_b_12_62432),
    .O(seg_15_18_local_g2_4_62592)
  );
  Span4Mux_v4 t1693 (
    .I(seg_16_19_sp4_h_l_36_51299),
    .O(seg_15_18_sp4_r_v_b_12_62432)
  );
  Span4Mux_h4 t1694 (
    .I(seg_12_19_sp4_h_l_47_35976),
    .O(seg_16_19_sp4_h_l_36_51299)
  );
  LocalMux t1695 (
    .I(seg_13_19_sp4_h_r_41_43642),
    .O(seg_13_19_local_g2_1_55052)
  );
  LocalMux t1696 (
    .I(seg_16_19_sp4_h_r_33_58970),
    .O(seg_16_19_local_g2_1_66543)
  );
  Span4Mux_h4 t1697 (
    .I(seg_14_19_sp4_h_l_43_43644),
    .O(seg_16_19_sp4_h_r_33_58970)
  );
  LocalMux t1698 (
    .I(seg_17_19_sp4_h_r_44_58970),
    .O(seg_17_19_local_g3_4_70385)
  );
  Span4Mux_h4 t1699 (
    .I(seg_14_19_sp4_h_l_43_43644),
    .O(seg_17_19_sp4_h_r_44_58970)
  );
  CascadeMux t17 (
    .I(net_16659),
    .O(net_16659_cascademuxed)
  );
  CascadeMux t170 (
    .I(net_43331),
    .O(net_43331_cascademuxed)
  );
  LocalMux t1700 (
    .I(seg_12_19_sp4_h_r_32_43646),
    .O(seg_12_19_local_g3_0_51228)
  );
  LocalMux t1701 (
    .I(seg_13_20_sp4_h_r_32_47600),
    .O(seg_13_20_local_g3_0_55182)
  );
  Span4Mux_h4 t1702 (
    .I(seg_11_20_sp4_v_b_8_43411),
    .O(seg_13_20_sp4_h_r_32_47600)
  );
  LocalMux t1703 (
    .I(seg_14_20_sp4_h_r_45_47600),
    .O(seg_14_20_local_g3_5_59017)
  );
  Span4Mux_h4 t1704 (
    .I(seg_11_20_sp4_v_b_8_43411),
    .O(seg_14_20_sp4_h_r_45_47600)
  );
  LocalMux t1705 (
    .I(seg_16_20_sp4_h_r_19_62920),
    .O(seg_16_20_local_g0_3_66652)
  );
  Span4Mux_h4 t1706 (
    .I(seg_15_20_sp4_h_l_47_47592),
    .O(seg_16_20_sp4_h_r_19_62920)
  );
  Span4Mux_h4 t1707 (
    .I(seg_11_20_sp4_v_b_10_43413),
    .O(seg_15_20_sp4_h_l_47_47592)
  );
  LocalMux t1708 (
    .I(seg_17_20_sp4_h_r_25_62913),
    .O(seg_17_20_local_g2_1_70497)
  );
  Span4Mux_h4 t1709 (
    .I(seg_15_20_sp4_h_l_47_47592),
    .O(seg_17_20_sp4_h_r_25_62913)
  );
  CascadeMux t171 (
    .I(net_43349),
    .O(net_43349_cascademuxed)
  );
  LocalMux t1710 (
    .I(seg_10_20_lutff_0_out_39793),
    .O(seg_10_20_local_g1_0_43673)
  );
  LocalMux t1711 (
    .I(seg_10_20_lutff_1_out_39794),
    .O(seg_10_20_local_g0_1_43666)
  );
  LocalMux t1712 (
    .I(seg_11_20_neigh_op_lft_1_39794),
    .O(seg_11_20_local_g1_1_47505)
  );
  LocalMux t1713 (
    .I(seg_10_20_lutff_2_out_39795),
    .O(seg_10_20_local_g3_2_43691)
  );
  LocalMux t1714 (
    .I(seg_11_20_neigh_op_lft_2_39795),
    .O(seg_11_20_local_g0_2_47498)
  );
  LocalMux t1715 (
    .I(seg_10_20_lutff_3_out_39796),
    .O(seg_10_20_local_g0_3_43668)
  );
  LocalMux t1716 (
    .I(seg_5_20_sp12_h_r_3_21400),
    .O(seg_5_20_local_g1_3_25152)
  );
  LocalMux t1717 (
    .I(seg_13_18_sp4_r_v_b_24_54896),
    .O(seg_13_18_local_g0_0_54912)
  );
  Span4Mux_v4 t1718 (
    .I(seg_14_20_sp4_h_l_37_43759),
    .O(seg_13_18_sp4_r_v_b_24_54896)
  );
  LocalMux t1719 (
    .I(seg_13_20_sp4_h_r_37_43759),
    .O(seg_13_20_local_g3_5_55187)
  );
  CascadeMux t172 (
    .I(net_43355),
    .O(net_43355_cascademuxed)
  );
  LocalMux t1720 (
    .I(seg_14_18_sp4_v_b_24_54896),
    .O(seg_14_18_local_g2_0_58758)
  );
  Span4Mux_v4 t1721 (
    .I(seg_14_20_sp4_h_l_37_43759),
    .O(seg_14_18_sp4_v_b_24_54896)
  );
  LocalMux t1722 (
    .I(seg_14_21_sp4_v_b_37_55388),
    .O(seg_14_21_local_g3_5_59140)
  );
  Span4Mux_v4 t1723 (
    .I(seg_14_20_sp4_h_l_37_43759),
    .O(seg_14_21_sp4_v_b_37_55388)
  );
  LocalMux t1724 (
    .I(seg_13_19_sp4_r_v_b_21_54904),
    .O(seg_13_19_local_g3_5_55064)
  );
  Span4Mux_v4 t1725 (
    .I(seg_14_20_sp4_h_l_39_43763),
    .O(seg_13_19_sp4_r_v_b_21_54904)
  );
  LocalMux t1726 (
    .I(seg_13_20_sp4_h_r_39_43763),
    .O(seg_13_20_local_g2_7_55181)
  );
  LocalMux t1727 (
    .I(seg_14_20_sp4_h_r_5_59089),
    .O(seg_14_20_local_g0_5_58993)
  );
  Span4Mux_h4 t1728 (
    .I(seg_14_20_sp4_h_l_39_43763),
    .O(seg_14_20_sp4_h_r_5_59089)
  );
  LocalMux t1729 (
    .I(seg_16_21_sp4_r_v_b_41_66883),
    .O(seg_16_21_local_g3_1_66797)
  );
  CascadeMux t173 (
    .I(net_43367),
    .O(net_43367_cascademuxed)
  );
  Span4Mux_v4 t1730 (
    .I(seg_17_20_sp4_h_l_46_55255),
    .O(seg_16_21_sp4_r_v_b_41_66883)
  );
  Span4Mux_h4 t1731 (
    .I(seg_13_20_sp4_h_l_46_39931),
    .O(seg_17_20_sp4_h_l_46_55255)
  );
  LocalMux t1732 (
    .I(seg_17_21_sp4_v_b_41_66883),
    .O(seg_17_21_local_g2_1_70620)
  );
  Span4Mux_v4 t1733 (
    .I(seg_17_20_sp4_h_l_46_55255),
    .O(seg_17_21_sp4_v_b_41_66883)
  );
  LocalMux t1734 (
    .I(seg_13_20_sp4_h_r_41_43765),
    .O(seg_13_20_local_g3_1_55183)
  );
  LocalMux t1735 (
    .I(seg_14_20_sp4_h_r_0_59082),
    .O(seg_14_20_local_g0_0_58988)
  );
  Span4Mux_h4 t1736 (
    .I(seg_14_20_sp4_h_l_41_43765),
    .O(seg_14_20_sp4_h_r_0_59082)
  );
  LocalMux t1737 (
    .I(seg_16_20_sp4_h_r_26_59086),
    .O(seg_16_20_local_g2_2_66667)
  );
  Span4Mux_h4 t1738 (
    .I(seg_14_20_sp4_h_l_43_43767),
    .O(seg_16_20_sp4_h_r_26_59086)
  );
  LocalMux t1739 (
    .I(seg_17_20_sp4_h_r_39_59086),
    .O(seg_17_20_local_g2_7_70503)
  );
  CascadeMux t174 (
    .I(net_43460),
    .O(net_43460_cascademuxed)
  );
  Span4Mux_h4 t1740 (
    .I(seg_14_20_sp4_h_l_43_43767),
    .O(seg_17_20_sp4_h_r_39_59086)
  );
  LocalMux t1741 (
    .I(seg_10_26_lutff_7_out_40538),
    .O(seg_10_26_local_g3_7_44434)
  );
  LocalMux t1742 (
    .I(seg_10_30_sp12_v_b_12_44250),
    .O(seg_10_30_local_g3_4_44923)
  );
  LocalMux t1743 (
    .I(seg_9_27_neigh_op_rgt_2_40656),
    .O(seg_9_27_local_g3_2_40721)
  );
  LocalMux t1744 (
    .I(seg_10_27_lutff_3_out_40657),
    .O(seg_10_27_local_g1_3_44537)
  );
  LocalMux t1745 (
    .I(seg_10_28_neigh_op_bot_4_40658),
    .O(seg_10_28_local_g0_4_44653)
  );
  LocalMux t1746 (
    .I(seg_10_27_lutff_5_out_40659),
    .O(seg_10_27_local_g1_5_44539)
  );
  LocalMux t1747 (
    .I(seg_10_27_lutff_6_out_40660),
    .O(seg_10_27_local_g0_6_44532)
  );
  LocalMux t1748 (
    .I(seg_10_28_neigh_op_bot_6_40660),
    .O(seg_10_28_local_g0_6_44655)
  );
  LocalMux t1749 (
    .I(seg_9_28_neigh_op_bnr_7_40661),
    .O(seg_9_28_local_g0_7_40825)
  );
  CascadeMux t175 (
    .I(net_43466),
    .O(net_43466_cascademuxed)
  );
  LocalMux t1750 (
    .I(seg_10_27_lutff_7_out_40661),
    .O(seg_10_27_local_g2_7_44549)
  );
  LocalMux t1751 (
    .I(seg_10_28_neigh_op_bot_7_40661),
    .O(seg_10_28_local_g0_7_44656)
  );
  LocalMux t1752 (
    .I(seg_10_28_lutff_2_out_40779),
    .O(seg_10_28_local_g3_2_44675)
  );
  LocalMux t1753 (
    .I(seg_9_28_neigh_op_rgt_3_40780),
    .O(seg_9_28_local_g2_3_40837)
  );
  LocalMux t1754 (
    .I(seg_10_27_neigh_op_top_3_40780),
    .O(seg_10_27_local_g0_3_44529)
  );
  LocalMux t1755 (
    .I(seg_10_28_lutff_3_out_40780),
    .O(seg_10_28_local_g1_3_44660)
  );
  LocalMux t1756 (
    .I(seg_10_27_neigh_op_top_7_40784),
    .O(seg_10_27_local_g0_7_44533)
  );
  LocalMux t1757 (
    .I(seg_10_28_lutff_7_out_40784),
    .O(seg_10_28_local_g1_7_44664)
  );
  LocalMux t1758 (
    .I(seg_10_30_sp4_v_b_2_40804),
    .O(seg_10_30_local_g1_2_44905)
  );
  LocalMux t1759 (
    .I(seg_9_29_neigh_op_rgt_0_40900),
    .O(seg_9_29_local_g2_0_40957)
  );
  CascadeMux t176 (
    .I(net_43484),
    .O(net_43484_cascademuxed)
  );
  LocalMux t1760 (
    .I(seg_9_29_neigh_op_rgt_0_40900),
    .O(seg_9_29_local_g3_0_40965)
  );
  LocalMux t1761 (
    .I(seg_9_30_neigh_op_bnr_0_40900),
    .O(seg_9_30_local_g1_0_41072)
  );
  LocalMux t1762 (
    .I(seg_10_29_lutff_0_out_40900),
    .O(seg_10_29_local_g2_0_44788)
  );
  LocalMux t1763 (
    .I(seg_10_30_neigh_op_bot_0_40900),
    .O(seg_10_30_local_g1_0_44903)
  );
  LocalMux t1764 (
    .I(seg_11_30_neigh_op_bnl_0_40900),
    .O(seg_11_30_local_g2_0_48742)
  );
  LocalMux t1765 (
    .I(seg_10_29_lutff_2_out_40902),
    .O(seg_10_29_local_g0_2_44774)
  );
  LocalMux t1766 (
    .I(seg_10_30_neigh_op_bot_2_40902),
    .O(seg_10_30_local_g0_2_44897)
  );
  LocalMux t1767 (
    .I(seg_11_29_neigh_op_lft_3_40903),
    .O(seg_11_29_local_g0_3_48606)
  );
  LocalMux t1768 (
    .I(seg_9_29_neigh_op_rgt_5_40905),
    .O(seg_9_29_local_g2_5_40962)
  );
  LocalMux t1769 (
    .I(seg_9_29_neigh_op_rgt_5_40905),
    .O(seg_9_29_local_g3_5_40970)
  );
  CascadeMux t177 (
    .I(net_43490),
    .O(net_43490_cascademuxed)
  );
  LocalMux t1770 (
    .I(seg_9_30_neigh_op_bnr_5_40905),
    .O(seg_9_30_local_g1_5_41077)
  );
  LocalMux t1771 (
    .I(seg_10_29_lutff_5_out_40905),
    .O(seg_10_29_local_g2_5_44793)
  );
  LocalMux t1772 (
    .I(seg_10_30_neigh_op_bot_5_40905),
    .O(seg_10_30_local_g1_5_44908)
  );
  LocalMux t1773 (
    .I(seg_11_29_neigh_op_lft_5_40905),
    .O(seg_11_29_local_g1_5_48616)
  );
  LocalMux t1774 (
    .I(seg_11_30_neigh_op_bnl_5_40905),
    .O(seg_11_30_local_g2_5_48747)
  );
  LocalMux t1775 (
    .I(seg_10_28_neigh_op_top_6_40906),
    .O(seg_10_28_local_g1_6_44663)
  );
  LocalMux t1776 (
    .I(seg_10_29_lutff_7_out_40907),
    .O(seg_10_29_local_g3_7_44803)
  );
  LocalMux t1777 (
    .I(seg_9_27_sp4_r_v_b_36_40801),
    .O(seg_9_27_local_g2_4_40715)
  );
  LocalMux t1778 (
    .I(seg_10_27_sp4_v_b_36_40801),
    .O(seg_10_27_local_g3_4_44554)
  );
  LocalMux t1779 (
    .I(seg_10_30_lutff_0_out_41023),
    .O(seg_10_30_local_g2_0_44911)
  );
  CascadeMux t178 (
    .I(net_43589),
    .O(net_43589_cascademuxed)
  );
  LocalMux t1780 (
    .I(seg_10_30_lutff_2_out_41025),
    .O(seg_10_30_local_g2_2_44913)
  );
  LocalMux t1781 (
    .I(seg_9_29_neigh_op_tnr_3_41026),
    .O(seg_9_29_local_g2_3_40960)
  );
  LocalMux t1782 (
    .I(seg_9_30_neigh_op_rgt_3_41026),
    .O(seg_9_30_local_g2_3_41083)
  );
  LocalMux t1783 (
    .I(seg_10_29_neigh_op_top_3_41026),
    .O(seg_10_29_local_g1_3_44783)
  );
  LocalMux t1784 (
    .I(seg_10_30_lutff_3_out_41026),
    .O(seg_10_30_local_g3_3_44922)
  );
  LocalMux t1785 (
    .I(seg_11_30_neigh_op_lft_3_41026),
    .O(seg_11_30_local_g1_3_48737)
  );
  LocalMux t1786 (
    .I(seg_9_29_neigh_op_tnr_4_41027),
    .O(seg_9_29_local_g2_4_40961)
  );
  LocalMux t1787 (
    .I(seg_9_30_neigh_op_rgt_4_41027),
    .O(seg_9_30_local_g2_4_41084)
  );
  LocalMux t1788 (
    .I(seg_10_29_neigh_op_top_4_41027),
    .O(seg_10_29_local_g1_4_44784)
  );
  LocalMux t1789 (
    .I(seg_10_30_lutff_4_out_41027),
    .O(seg_10_30_local_g0_4_44899)
  );
  CascadeMux t179 (
    .I(net_43613),
    .O(net_43613_cascademuxed)
  );
  LocalMux t1790 (
    .I(seg_10_30_lutff_4_out_41027),
    .O(seg_10_30_local_g1_4_44907)
  );
  LocalMux t1791 (
    .I(seg_11_30_neigh_op_lft_4_41027),
    .O(seg_11_30_local_g1_4_48738)
  );
  LocalMux t1792 (
    .I(seg_10_30_lutff_6_out_41029),
    .O(seg_10_30_local_g2_6_44917)
  );
  LocalMux t1793 (
    .I(seg_10_30_lutff_7_out_41030),
    .O(seg_10_30_local_g3_7_44926)
  );
  LocalMux t1794 (
    .I(seg_10_8_neigh_op_bnr_0_42025),
    .O(seg_10_8_local_g1_0_42197)
  );
  LocalMux t1795 (
    .I(seg_11_7_lutff_0_out_42025),
    .O(seg_11_7_local_g3_0_45921)
  );
  LocalMux t1796 (
    .I(seg_11_8_neigh_op_bot_0_42025),
    .O(seg_11_8_local_g1_0_46028)
  );
  LocalMux t1797 (
    .I(seg_12_8_neigh_op_bnl_0_42025),
    .O(seg_12_8_local_g3_0_49875)
  );
  LocalMux t1798 (
    .I(seg_11_7_lutff_2_out_42027),
    .O(seg_11_7_local_g1_2_45907)
  );
  LocalMux t1799 (
    .I(seg_11_7_lutff_7_out_42032),
    .O(seg_11_7_local_g1_7_45912)
  );
  CascadeMux t18 (
    .I(net_16665),
    .O(net_16665_cascademuxed)
  );
  CascadeMux t180 (
    .I(net_43619),
    .O(net_43619_cascademuxed)
  );
  LocalMux t1800 (
    .I(seg_9_8_sp4_h_r_17_34627),
    .O(seg_9_8_local_g1_1_38367)
  );
  Span4Mux_h4 t1801 (
    .I(seg_12_8_sp4_v_b_4_45762),
    .O(seg_9_8_sp4_h_r_17_34627)
  );
  LocalMux t1802 (
    .I(seg_11_9_neigh_op_bot_2_42150),
    .O(seg_11_9_local_g0_2_46145)
  );
  LocalMux t1803 (
    .I(seg_11_9_neigh_op_bot_3_42151),
    .O(seg_11_9_local_g0_3_46146)
  );
  LocalMux t1804 (
    .I(seg_11_9_neigh_op_bot_4_42152),
    .O(seg_11_9_local_g0_4_46147)
  );
  LocalMux t1805 (
    .I(seg_10_8_neigh_op_rgt_5_42153),
    .O(seg_10_8_local_g2_5_42210)
  );
  LocalMux t1806 (
    .I(seg_10_8_neigh_op_rgt_6_42154),
    .O(seg_10_8_local_g2_6_42211)
  );
  LocalMux t1807 (
    .I(seg_10_8_neigh_op_rgt_7_42155),
    .O(seg_10_8_local_g3_7_42220)
  );
  LocalMux t1808 (
    .I(seg_11_8_neigh_op_top_0_42271),
    .O(seg_11_8_local_g0_0_46020)
  );
  LocalMux t1809 (
    .I(seg_11_8_neigh_op_top_1_42272),
    .O(seg_11_8_local_g0_1_46021)
  );
  CascadeMux t181 (
    .I(net_43706),
    .O(net_43706_cascademuxed)
  );
  LocalMux t1810 (
    .I(seg_11_8_neigh_op_top_3_42274),
    .O(seg_11_8_local_g0_3_46023)
  );
  LocalMux t1811 (
    .I(seg_11_9_lutff_4_out_42275),
    .O(seg_11_9_local_g1_4_46155)
  );
  LocalMux t1812 (
    .I(seg_11_9_lutff_5_out_42276),
    .O(seg_11_9_local_g1_5_46156)
  );
  LocalMux t1813 (
    .I(seg_11_9_lutff_6_out_42277),
    .O(seg_11_9_local_g2_6_46165)
  );
  LocalMux t1814 (
    .I(seg_11_10_neigh_op_bot_7_42278),
    .O(seg_11_10_local_g0_7_46273)
  );
  LocalMux t1815 (
    .I(seg_9_8_sp4_r_v_b_16_38222),
    .O(seg_9_8_local_g3_0_38382)
  );
  Span4Mux_v4 t1816 (
    .I(seg_10_9_sp4_h_r_5_42413),
    .O(seg_9_8_sp4_r_v_b_16_38222)
  );
  LocalMux t1817 (
    .I(seg_9_8_sp4_r_v_b_17_38223),
    .O(seg_9_8_local_g3_1_38383)
  );
  Span4Mux_v4 t1818 (
    .I(seg_10_9_sp4_h_r_11_42409),
    .O(seg_9_8_sp4_r_v_b_17_38223)
  );
  LocalMux t1819 (
    .I(seg_9_8_sp4_v_b_14_34389),
    .O(seg_9_8_local_g0_6_38364)
  );
  CascadeMux t182 (
    .I(net_43718),
    .O(net_43718_cascademuxed)
  );
  Span4Mux_v4 t1820 (
    .I(seg_9_9_sp4_h_r_10_38577),
    .O(seg_9_8_sp4_v_b_14_34389)
  );
  LocalMux t1821 (
    .I(seg_12_11_neigh_op_bnl_4_42398),
    .O(seg_12_11_local_g2_4_50240)
  );
  LocalMux t1822 (
    .I(seg_11_10_lutff_5_out_42399),
    .O(seg_11_10_local_g1_5_46279)
  );
  LocalMux t1823 (
    .I(seg_11_9_neigh_op_top_6_42400),
    .O(seg_11_9_local_g0_6_46149)
  );
  LocalMux t1824 (
    .I(seg_11_10_lutff_7_out_42401),
    .O(seg_11_10_local_g3_7_46297)
  );
  LocalMux t1825 (
    .I(seg_13_9_sp4_r_v_b_18_53671),
    .O(seg_13_9_local_g3_2_53831)
  );
  Span4Mux_v4 t1826 (
    .I(seg_14_10_sp4_h_l_36_42530),
    .O(seg_13_9_sp4_r_v_b_18_53671)
  );
  LocalMux t1827 (
    .I(seg_14_8_sp4_v_b_31_53671),
    .O(seg_14_8_local_g2_7_57535)
  );
  Span4Mux_v4 t1828 (
    .I(seg_14_10_sp4_h_l_36_42530),
    .O(seg_14_8_sp4_v_b_31_53671)
  );
  LocalMux t1829 (
    .I(seg_14_8_sp4_v_b_31_53671),
    .O(seg_14_8_local_g3_7_57543)
  );
  CascadeMux t183 (
    .I(net_44561),
    .O(net_44561_cascademuxed)
  );
  LocalMux t1830 (
    .I(seg_15_10_sp4_h_r_19_57860),
    .O(seg_15_10_local_g0_3_61591)
  );
  Span4Mux_h4 t1831 (
    .I(seg_14_10_sp4_h_l_38_42534),
    .O(seg_15_10_sp4_h_r_19_57860)
  );
  LocalMux t1832 (
    .I(seg_13_12_sp4_v_b_24_50327),
    .O(seg_13_12_local_g2_0_54190)
  );
  Span4Mux_v4 t1833 (
    .I(seg_13_10_sp4_h_l_37_38698),
    .O(seg_13_12_sp4_v_b_24_50327)
  );
  LocalMux t1834 (
    .I(seg_13_14_sp4_v_b_0_50327),
    .O(seg_13_14_local_g1_0_54428)
  );
  Span4Mux_v4 t1835 (
    .I(seg_13_10_sp4_h_l_37_38698),
    .O(seg_13_14_sp4_v_b_0_50327)
  );
  LocalMux t1836 (
    .I(seg_13_19_sp4_v_b_43_51317),
    .O(seg_13_19_local_g3_3_55062)
  );
  Span4Mux_v4 t1837 (
    .I(seg_13_18_sp4_v_b_3_50820),
    .O(seg_13_19_sp4_v_b_43_51317)
  );
  Span4Mux_v4 t1838 (
    .I(seg_13_14_sp4_v_b_0_50327),
    .O(seg_13_18_sp4_v_b_3_50820)
  );
  LocalMux t1839 (
    .I(seg_11_14_sp4_v_b_2_42667),
    .O(seg_11_14_local_g1_2_46768)
  );
  CascadeMux t184 (
    .I(net_44567),
    .O(net_44567_cascademuxed)
  );
  Span4Mux_v4 t1840 (
    .I(seg_11_10_sp4_h_r_8_46370),
    .O(seg_11_14_sp4_v_b_2_42667)
  );
  LocalMux t1841 (
    .I(seg_11_18_sp4_v_b_10_43167),
    .O(seg_11_18_local_g0_2_47252)
  );
  Span4Mux_v4 t1842 (
    .I(seg_11_14_sp4_v_b_2_42667),
    .O(seg_11_18_sp4_v_b_10_43167)
  );
  LocalMux t1843 (
    .I(seg_14_10_sp4_h_r_45_46370),
    .O(seg_14_10_local_g2_5_57779)
  );
  LocalMux t1844 (
    .I(seg_14_13_sp4_r_v_b_21_57996),
    .O(seg_14_13_local_g3_5_58156)
  );
  Span4Mux_v4 t1845 (
    .I(seg_15_10_sp4_h_l_45_46370),
    .O(seg_14_13_sp4_r_v_b_21_57996)
  );
  LocalMux t1846 (
    .I(seg_15_10_sp4_h_r_4_61688),
    .O(seg_15_10_local_g1_4_61600)
  );
  Span4Mux_h4 t1847 (
    .I(seg_15_10_sp4_h_l_45_46370),
    .O(seg_15_10_sp4_h_r_4_61688)
  );
  LocalMux t1848 (
    .I(seg_15_16_sp4_v_b_28_58484),
    .O(seg_15_16_local_g2_4_62346)
  );
  Span4Mux_v4 t1849 (
    .I(seg_15_14_sp4_v_b_8_57996),
    .O(seg_15_16_sp4_v_b_28_58484)
  );
  CascadeMux t185 (
    .I(net_44579),
    .O(net_44579_cascademuxed)
  );
  Span4Mux_v4 t1850 (
    .I(seg_15_10_sp4_h_l_45_46370),
    .O(seg_15_14_sp4_v_b_8_57996)
  );
  LocalMux t1851 (
    .I(seg_15_17_sp4_v_b_17_58484),
    .O(seg_15_17_local_g1_1_62458)
  );
  Span4Mux_v4 t1852 (
    .I(seg_15_14_sp4_v_b_8_57996),
    .O(seg_15_17_sp4_v_b_17_58484)
  );
  LocalMux t1853 (
    .I(seg_15_18_sp4_v_b_4_58484),
    .O(seg_15_18_local_g1_4_62584)
  );
  Span4Mux_v4 t1854 (
    .I(seg_15_14_sp4_v_b_8_57996),
    .O(seg_15_18_sp4_v_b_4_58484)
  );
  LocalMux t1855 (
    .I(seg_10_7_sp4_h_r_24_34498),
    .O(seg_10_7_local_g2_0_42082)
  );
  Span4Mux_h4 t1856 (
    .I(seg_12_7_sp4_v_t_37_46127),
    .O(seg_10_7_sp4_h_r_24_34498)
  );
  LocalMux t1857 (
    .I(seg_12_8_sp4_v_b_37_46127),
    .O(seg_12_8_local_g3_5_49880)
  );
  LocalMux t1858 (
    .I(seg_14_7_sp4_h_r_29_49829),
    .O(seg_14_7_local_g2_5_57410)
  );
  Span4Mux_h4 t1859 (
    .I(seg_12_7_sp4_v_t_37_46127),
    .O(seg_14_7_sp4_h_r_29_49829)
  );
  CascadeMux t186 (
    .I(net_44696),
    .O(net_44696_cascademuxed)
  );
  LocalMux t1860 (
    .I(seg_11_19_sp4_r_v_b_16_47237),
    .O(seg_11_19_local_g3_0_47397)
  );
  Span4Mux_v4 t1861 (
    .I(seg_12_16_sp4_v_b_9_46749),
    .O(seg_11_19_sp4_r_v_b_16_47237)
  );
  Span4Mux_v4 t1862 (
    .I(seg_12_12_sp4_v_b_1_46249),
    .O(seg_12_16_sp4_v_b_9_46749)
  );
  LocalMux t1863 (
    .I(seg_12_15_sp4_v_b_17_46746),
    .O(seg_12_15_local_g0_1_50713)
  );
  Span4Mux_v4 t1864 (
    .I(seg_12_12_sp4_v_b_1_46249),
    .O(seg_12_15_sp4_v_b_17_46746)
  );
  LocalMux t1865 (
    .I(seg_12_15_sp4_v_b_20_46749),
    .O(seg_12_15_local_g0_4_50716)
  );
  Span4Mux_v4 t1866 (
    .I(seg_12_12_sp4_v_b_1_46249),
    .O(seg_12_15_sp4_v_b_20_46749)
  );
  LocalMux t1867 (
    .I(seg_13_20_sp4_h_r_22_51424),
    .O(seg_13_20_local_g1_6_55172)
  );
  Span4Mux_h4 t1868 (
    .I(seg_12_20_sp4_v_b_5_47237),
    .O(seg_13_20_sp4_h_r_22_51424)
  );
  Span4Mux_v4 t1869 (
    .I(seg_12_16_sp4_v_b_9_46749),
    .O(seg_12_20_sp4_v_b_5_47237)
  );
  CascadeMux t187 (
    .I(net_44702),
    .O(net_44702_cascademuxed)
  );
  LocalMux t1870 (
    .I(seg_15_19_sp4_r_v_b_20_62563),
    .O(seg_15_19_local_g3_4_62723)
  );
  Span4Mux_v4 t1871 (
    .I(seg_16_16_sp4_v_b_1_62063),
    .O(seg_15_19_sp4_r_v_b_20_62563)
  );
  Span4Mux_v4 t1872 (
    .I(seg_16_12_sp4_h_l_36_50438),
    .O(seg_16_16_sp4_v_b_1_62063)
  );
  Span4Mux_h4 t1873 (
    .I(seg_12_12_sp4_v_b_1_46249),
    .O(seg_16_12_sp4_h_l_36_50438)
  );
  LocalMux t1874 (
    .I(seg_16_16_sp4_v_b_1_62063),
    .O(seg_16_16_local_g0_1_66158)
  );
  LocalMux t1875 (
    .I(seg_16_19_sp4_v_b_20_62563),
    .O(seg_16_19_local_g1_4_66538)
  );
  Span4Mux_v4 t1876 (
    .I(seg_16_16_sp4_v_b_1_62063),
    .O(seg_16_19_sp4_v_b_20_62563)
  );
  LocalMux t1877 (
    .I(seg_16_20_sp4_v_b_9_62563),
    .O(seg_16_20_local_g1_1_66658)
  );
  Span4Mux_v4 t1878 (
    .I(seg_16_16_sp4_v_b_1_62063),
    .O(seg_16_20_sp4_v_b_9_62563)
  );
  LocalMux t1879 (
    .I(seg_20_16_sp4_v_b_5_77117),
    .O(seg_20_16_local_g0_5_80855)
  );
  CascadeMux t188 (
    .I(net_44714),
    .O(net_44714_cascademuxed)
  );
  Span4Mux_v4 t1880 (
    .I(seg_20_12_sp4_h_l_40_65766),
    .O(seg_20_16_sp4_v_b_5_77117)
  );
  Span4Mux_h4 t1881 (
    .I(seg_16_12_sp4_h_l_40_50444),
    .O(seg_20_12_sp4_h_l_40_65766)
  );
  Span4Mux_h4 t1882 (
    .I(seg_12_12_sp4_v_b_5_46253),
    .O(seg_16_12_sp4_h_l_40_50444)
  );
  LocalMux t1883 (
    .I(seg_15_20_sp4_r_v_b_7_62561),
    .O(seg_15_20_local_g1_7_62833)
  );
  Span4Mux_v4 t1884 (
    .I(seg_16_16_sp4_v_b_7_62069),
    .O(seg_15_20_sp4_r_v_b_7_62561)
  );
  Span4Mux_v4 t1885 (
    .I(seg_16_12_sp4_h_l_42_50446),
    .O(seg_16_16_sp4_v_b_7_62069)
  );
  Span4Mux_h4 t1886 (
    .I(seg_12_12_sp4_v_b_7_46255),
    .O(seg_16_12_sp4_h_l_42_50446)
  );
  LocalMux t1887 (
    .I(seg_11_10_sp4_r_v_b_33_46257),
    .O(seg_11_10_local_g0_2_46268)
  );
  GlobalMux t1888 (
    .I(seg_13_31_local_g1_4_56536_i3),
    .O(seg_9_11_glb_netwk_1_6)
  );
  gio2CtrlBuf t1889 (
    .I(seg_13_31_local_g1_4_56536_i2),
    .O(seg_13_31_local_g1_4_56536_i3)
  );
  CascadeMux t189 (
    .I(net_44726),
    .O(net_44726_cascademuxed)
  );
  ICE_GB t1890 (
    .GLOBALBUFFEROUTPUT(seg_13_31_local_g1_4_56536_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_13_31_local_g1_4_56536_i1)
  );
  IoInMux t1891 (
    .I(seg_13_31_local_g1_4_56536),
    .O(seg_13_31_local_g1_4_56536_i1)
  );
  LocalMux t1892 (
    .I(seg_13_31_span4_horz_r_4_52709),
    .O(seg_13_31_local_g1_4_56536)
  );
  IoSpan4Mux t1893 (
    .I(seg_12_31_span4_vert_25_48828),
    .O(seg_13_31_span4_horz_r_4_52709)
  );
  Span4Mux_v4 t1894 (
    .I(seg_12_29_sp4_v_b_1_48340),
    .O(seg_12_31_span4_vert_25_48828)
  );
  Span4Mux_v4 t1895 (
    .I(seg_12_25_sp4_v_b_1_47848),
    .O(seg_12_29_sp4_v_b_1_48340)
  );
  Span4Mux_v4 t1896 (
    .I(seg_12_21_sp4_v_b_1_47356),
    .O(seg_12_25_sp4_v_b_1_47848)
  );
  Span4Mux_v4 t1897 (
    .I(seg_12_17_sp4_v_b_5_46868),
    .O(seg_12_21_sp4_v_b_1_47356)
  );
  Span4Mux_v4 t1898 (
    .I(seg_12_13_sp4_v_b_2_46375),
    .O(seg_12_17_sp4_v_b_5_46868)
  );
  LocalMux t1899 (
    .I(seg_11_12_sp4_r_v_b_17_46377),
    .O(seg_11_12_local_g3_1_46537)
  );
  CascadeMux t19 (
    .I(net_16689),
    .O(net_16689_cascademuxed)
  );
  CascadeMux t190 (
    .I(net_44807),
    .O(net_44807_cascademuxed)
  );
  LocalMux t1900 (
    .I(seg_13_13_sp4_h_r_23_50562),
    .O(seg_13_13_local_g1_7_54312)
  );
  Span4Mux_h4 t1901 (
    .I(seg_12_13_sp4_v_b_4_46377),
    .O(seg_13_13_sp4_h_r_23_50562)
  );
  LocalMux t1902 (
    .I(seg_12_21_sp4_v_b_10_47367),
    .O(seg_12_21_local_g0_2_51452)
  );
  Span4Mux_v4 t1903 (
    .I(seg_12_17_sp4_v_b_10_46875),
    .O(seg_12_21_sp4_v_b_10_47367)
  );
  Span4Mux_v4 t1904 (
    .I(seg_12_13_sp4_v_b_10_46383),
    .O(seg_12_17_sp4_v_b_10_46875)
  );
  LocalMux t1905 (
    .I(seg_12_14_sp4_v_b_9_46503),
    .O(seg_12_14_local_g1_1_50598)
  );
  Span4Mux_v4 t1906 (
    .I(seg_12_10_sp4_v_b_9_46011),
    .O(seg_12_14_sp4_v_b_9_46503)
  );
  LocalMux t1907 (
    .I(seg_12_18_sp4_v_b_9_46995),
    .O(seg_12_18_local_g0_1_51082)
  );
  Span4Mux_v4 t1908 (
    .I(seg_12_14_sp4_v_b_9_46503),
    .O(seg_12_18_sp4_v_b_9_46995)
  );
  LocalMux t1909 (
    .I(seg_13_14_sp4_h_r_14_50688),
    .O(seg_13_14_local_g1_6_54434)
  );
  CascadeMux t191 (
    .I(net_44825),
    .O(net_44825_cascademuxed)
  );
  Span4Mux_h4 t1910 (
    .I(seg_12_14_sp4_v_b_9_46503),
    .O(seg_13_14_sp4_h_r_14_50688)
  );
  LocalMux t1911 (
    .I(seg_10_8_sp4_r_v_b_36_42295),
    .O(seg_10_8_local_g2_4_42209)
  );
  LocalMux t1912 (
    .I(seg_11_7_sp4_h_r_6_45999),
    .O(seg_11_7_local_g1_6_45911)
  );
  Span4Mux_h4 t1913 (
    .I(seg_11_7_sp4_v_t_36_42295),
    .O(seg_11_7_sp4_h_r_6_45999)
  );
  LocalMux t1914 (
    .I(seg_14_15_sp4_r_v_b_16_58237),
    .O(seg_14_15_local_g3_0_58397)
  );
  Span4Mux_v4 t1915 (
    .I(seg_15_12_sp4_h_l_37_46606),
    .O(seg_14_15_sp4_r_v_b_16_58237)
  );
  Span4Mux_h4 t1916 (
    .I(seg_11_12_sp4_v_b_0_42419),
    .O(seg_15_12_sp4_h_l_37_46606)
  );
  LocalMux t1917 (
    .I(seg_14_16_sp4_r_v_b_5_58237),
    .O(seg_14_16_local_g1_5_58509)
  );
  Span4Mux_v4 t1918 (
    .I(seg_15_12_sp4_h_l_37_46606),
    .O(seg_14_16_sp4_r_v_b_5_58237)
  );
  LocalMux t1919 (
    .I(seg_14_19_sp4_r_v_b_21_58734),
    .O(seg_14_19_local_g3_5_58894)
  );
  CascadeMux t192 (
    .I(net_44837),
    .O(net_44837_cascademuxed)
  );
  Span4Mux_v4 t1920 (
    .I(seg_15_16_sp4_v_b_5_58237),
    .O(seg_14_19_sp4_r_v_b_21_58734)
  );
  Span4Mux_v4 t1921 (
    .I(seg_15_12_sp4_h_l_37_46606),
    .O(seg_15_16_sp4_v_b_5_58237)
  );
  LocalMux t1922 (
    .I(seg_14_20_sp4_r_v_b_8_58734),
    .O(seg_14_20_local_g2_0_59004)
  );
  Span4Mux_v4 t1923 (
    .I(seg_15_16_sp4_v_b_5_58237),
    .O(seg_14_20_sp4_r_v_b_8_58734)
  );
  LocalMux t1924 (
    .I(seg_11_13_sp4_v_b_5_42545),
    .O(seg_11_13_local_g0_5_46640)
  );
  LocalMux t1925 (
    .I(seg_18_16_sp4_r_v_b_22_73689),
    .O(seg_18_16_local_g3_6_73849)
  );
  Span4Mux_v4 t1926 (
    .I(seg_19_13_sp4_h_l_46_62054),
    .O(seg_18_16_sp4_r_v_b_22_73689)
  );
  Span4Mux_h4 t1927 (
    .I(seg_15_13_sp4_h_l_38_46734),
    .O(seg_19_13_sp4_h_l_46_62054)
  );
  Span4Mux_h4 t1928 (
    .I(seg_11_13_sp4_v_b_9_42549),
    .O(seg_15_13_sp4_h_l_38_46734)
  );
  LocalMux t1929 (
    .I(seg_10_11_neigh_op_rgt_2_42519),
    .O(seg_10_11_local_g2_2_42576)
  );
  CascadeMux t193 (
    .I(net_44843),
    .O(net_44843_cascademuxed)
  );
  LocalMux t1930 (
    .I(seg_12_11_neigh_op_lft_2_42519),
    .O(seg_12_11_local_g1_2_50230)
  );
  LocalMux t1931 (
    .I(seg_10_11_neigh_op_rgt_7_42524),
    .O(seg_10_11_local_g2_7_42581)
  );
  LocalMux t1932 (
    .I(seg_12_11_neigh_op_lft_7_42524),
    .O(seg_12_11_local_g0_7_50227)
  );
  LocalMux t1933 (
    .I(seg_11_12_lutff_2_out_42642),
    .O(seg_11_12_local_g0_2_46514)
  );
  LocalMux t1934 (
    .I(seg_10_12_neigh_op_rgt_6_42646),
    .O(seg_10_12_local_g2_6_42703)
  );
  LocalMux t1935 (
    .I(seg_11_13_neigh_op_bot_7_42647),
    .O(seg_11_13_local_g0_7_46642)
  );
  LocalMux t1936 (
    .I(seg_14_13_sp4_v_b_38_54405),
    .O(seg_14_13_local_g2_6_58149)
  );
  Span4Mux_v4 t1937 (
    .I(seg_14_12_sp4_h_l_38_42780),
    .O(seg_14_13_sp4_v_b_38_54405)
  );
  LocalMux t1938 (
    .I(seg_14_12_sp4_h_r_39_46610),
    .O(seg_14_12_local_g3_7_58035)
  );
  LocalMux t1939 (
    .I(seg_13_12_sp4_h_r_44_42786),
    .O(seg_13_12_local_g3_4_54202)
  );
  CascadeMux t194 (
    .I(net_44849),
    .O(net_44849_cascademuxed)
  );
  LocalMux t1940 (
    .I(seg_14_12_sp4_h_r_43_46614),
    .O(seg_14_12_local_g3_3_58031)
  );
  LocalMux t1941 (
    .I(seg_15_13_sp4_v_b_36_58233),
    .O(seg_15_13_local_g3_4_61985)
  );
  Span4Mux_v4 t1942 (
    .I(seg_15_12_sp4_h_l_45_46616),
    .O(seg_15_13_sp4_v_b_36_58233)
  );
  LocalMux t1943 (
    .I(seg_10_13_neigh_op_rgt_3_42766),
    .O(seg_10_13_local_g2_3_42823)
  );
  LocalMux t1944 (
    .I(seg_10_13_neigh_op_rgt_7_42770),
    .O(seg_10_13_local_g3_7_42835)
  );
  LocalMux t1945 (
    .I(seg_14_13_sp12_h_r_9_42895),
    .O(seg_14_13_local_g1_1_58136)
  );
  LocalMux t1946 (
    .I(seg_15_13_sp4_h_r_17_58227),
    .O(seg_15_13_local_g1_1_61966)
  );
  Span4Mux_h4 t1947 (
    .I(seg_14_13_sp4_h_l_36_42899),
    .O(seg_15_13_sp4_h_r_17_58227)
  );
  LocalMux t1948 (
    .I(seg_14_13_sp4_h_r_39_46733),
    .O(seg_14_13_local_g2_7_58150)
  );
  LocalMux t1949 (
    .I(seg_15_13_sp4_h_r_27_54396),
    .O(seg_15_13_local_g3_3_61984)
  );
  CascadeMux t195 (
    .I(net_44930),
    .O(net_44930_cascademuxed)
  );
  Span4Mux_h4 t1950 (
    .I(seg_13_13_sp4_h_l_37_39067),
    .O(seg_15_13_sp4_h_r_27_54396)
  );
  LocalMux t1951 (
    .I(seg_15_13_sp4_h_r_32_54401),
    .O(seg_15_13_local_g2_0_61973)
  );
  Span4Mux_h4 t1952 (
    .I(seg_13_13_sp4_h_l_45_39077),
    .O(seg_15_13_sp4_h_r_32_54401)
  );
  LocalMux t1953 (
    .I(seg_14_13_sp4_h_r_41_46735),
    .O(seg_14_13_local_g2_1_58144)
  );
  LocalMux t1954 (
    .I(seg_11_14_lutff_0_out_42886),
    .O(seg_11_14_local_g2_0_46774)
  );
  LocalMux t1955 (
    .I(seg_12_13_neigh_op_tnl_2_42888),
    .O(seg_12_13_local_g2_2_50484)
  );
  LocalMux t1956 (
    .I(seg_12_13_neigh_op_tnl_3_42889),
    .O(seg_12_13_local_g2_3_50485)
  );
  LocalMux t1957 (
    .I(seg_12_14_neigh_op_lft_4_42890),
    .O(seg_12_14_local_g1_4_50601)
  );
  LocalMux t1958 (
    .I(seg_11_14_lutff_6_out_42892),
    .O(seg_11_14_local_g2_6_46780)
  );
  LocalMux t1959 (
    .I(seg_14_14_sp4_h_r_6_58352),
    .O(seg_14_14_local_g1_6_58264)
  );
  CascadeMux t196 (
    .I(net_44942),
    .O(net_44942_cascademuxed)
  );
  Span4Mux_h4 t1960 (
    .I(seg_14_14_sp4_h_l_38_43026),
    .O(seg_14_14_sp4_h_r_6_58352)
  );
  LocalMux t1961 (
    .I(seg_14_14_sp4_h_r_39_46856),
    .O(seg_14_14_local_g2_7_58273)
  );
  LocalMux t1962 (
    .I(seg_16_15_sp4_v_b_14_62065),
    .O(seg_16_15_local_g0_6_66040)
  );
  Span4Mux_v4 t1963 (
    .I(seg_16_16_sp4_h_l_44_50940),
    .O(seg_16_15_sp4_v_b_14_62065)
  );
  Span4Mux_h4 t1964 (
    .I(seg_12_16_sp4_v_b_3_46743),
    .O(seg_16_16_sp4_h_l_44_50940)
  );
  LocalMux t1965 (
    .I(seg_12_15_neigh_op_lft_2_43011),
    .O(seg_12_15_local_g1_2_50722)
  );
  LocalMux t1966 (
    .I(seg_12_14_neigh_op_tnl_4_43013),
    .O(seg_12_14_local_g3_4_50617)
  );
  LocalMux t1967 (
    .I(seg_12_15_neigh_op_lft_4_43013),
    .O(seg_12_15_local_g1_4_50724)
  );
  LocalMux t1968 (
    .I(seg_12_15_neigh_op_lft_6_43015),
    .O(seg_12_15_local_g0_6_50718)
  );
  LocalMux t1969 (
    .I(seg_10_13_sp4_r_v_b_30_42794),
    .O(seg_10_13_local_g0_6_42810)
  );
  CascadeMux t197 (
    .I(net_44948),
    .O(net_44948_cascademuxed)
  );
  LocalMux t1970 (
    .I(seg_10_17_neigh_op_bnr_5_43137),
    .O(seg_10_17_local_g1_5_43309)
  );
  LocalMux t1971 (
    .I(seg_11_16_lutff_5_out_43137),
    .O(seg_11_16_local_g0_5_47009)
  );
  LocalMux t1972 (
    .I(seg_13_16_sp4_h_r_34_47100),
    .O(seg_13_16_local_g3_2_54692)
  );
  LocalMux t1973 (
    .I(seg_10_12_sp4_h_r_35_35116),
    .O(seg_10_12_local_g3_3_42708)
  );
  Span4Mux_h4 t1974 (
    .I(seg_12_12_sp4_v_t_46_46751),
    .O(seg_10_12_sp4_h_r_35_35116)
  );
  LocalMux t1975 (
    .I(seg_11_11_sp4_r_v_b_22_46259),
    .O(seg_11_11_local_g3_6_46419)
  );
  Span4Mux_v4 t1976 (
    .I(seg_12_12_sp4_v_t_46_46751),
    .O(seg_11_11_sp4_r_v_b_22_46259)
  );
  LocalMux t1977 (
    .I(seg_12_11_sp4_v_b_22_46259),
    .O(seg_12_11_local_g1_6_50234)
  );
  Span4Mux_v4 t1978 (
    .I(seg_12_12_sp4_v_t_46_46751),
    .O(seg_12_11_sp4_v_b_22_46259)
  );
  LocalMux t1979 (
    .I(seg_12_12_sp4_h_r_11_50440),
    .O(seg_12_12_local_g0_3_50346)
  );
  CascadeMux t198 (
    .I(net_44954),
    .O(net_44954_cascademuxed)
  );
  Span4Mux_h4 t1980 (
    .I(seg_12_12_sp4_v_t_46_46751),
    .O(seg_12_12_sp4_h_r_11_50440)
  );
  LocalMux t1981 (
    .I(seg_15_11_sp4_r_v_b_22_61581),
    .O(seg_15_11_local_g3_6_61741)
  );
  Span4Mux_v4 t1982 (
    .I(seg_16_12_sp4_h_l_46_50440),
    .O(seg_15_11_sp4_r_v_b_22_61581)
  );
  Span4Mux_h4 t1983 (
    .I(seg_12_12_sp4_v_t_46_46751),
    .O(seg_16_12_sp4_h_l_46_50440)
  );
  LocalMux t1984 (
    .I(seg_16_11_sp4_v_b_22_61581),
    .O(seg_16_11_local_g0_6_65548)
  );
  Span4Mux_v4 t1985 (
    .I(seg_16_12_sp4_h_l_46_50440),
    .O(seg_16_11_sp4_v_b_22_61581)
  );
  LocalMux t1986 (
    .I(seg_14_15_sp4_h_r_30_50814),
    .O(seg_14_15_local_g3_6_58403)
  );
  Span4Mux_h4 t1987 (
    .I(seg_12_15_sp4_v_t_43_47117),
    .O(seg_14_15_sp4_h_r_30_50814)
  );
  LocalMux t1988 (
    .I(seg_10_17_neigh_op_rgt_1_43256),
    .O(seg_10_17_local_g3_1_43321)
  );
  LocalMux t1989 (
    .I(seg_11_17_lutff_1_out_43256),
    .O(seg_11_17_local_g0_1_47128)
  );
  CascadeMux t199 (
    .I(net_44966),
    .O(net_44966_cascademuxed)
  );
  LocalMux t1990 (
    .I(seg_13_16_sp4_r_v_b_12_54526),
    .O(seg_13_16_local_g2_4_54686)
  );
  Span4Mux_v4 t1991 (
    .I(seg_14_17_sp4_h_l_42_43399),
    .O(seg_13_16_sp4_r_v_b_12_54526)
  );
  LocalMux t1992 (
    .I(seg_11_16_sp4_v_b_18_43039),
    .O(seg_11_16_local_g0_2_47006)
  );
  Span4Mux_v4 t1993 (
    .I(seg_11_17_sp4_h_r_2_47225),
    .O(seg_11_16_sp4_v_b_18_43039)
  );
  LocalMux t1994 (
    .I(seg_12_12_sp4_v_b_42_46624),
    .O(seg_12_12_local_g2_2_50361)
  );
  Span4Mux_v4 t1995 (
    .I(seg_12_15_sp4_v_t_46_47120),
    .O(seg_12_12_sp4_v_b_42_46624)
  );
  LocalMux t1996 (
    .I(seg_13_11_sp4_h_r_13_50314),
    .O(seg_13_11_local_g1_5_54064)
  );
  Span4Mux_h4 t1997 (
    .I(seg_12_11_sp4_v_t_42_46624),
    .O(seg_13_11_sp4_h_r_13_50314)
  );
  Span4Mux_v4 t1998 (
    .I(seg_12_15_sp4_v_t_46_47120),
    .O(seg_12_11_sp4_v_t_42_46624)
  );
  LocalMux t1999 (
    .I(seg_14_11_sp4_h_r_24_50314),
    .O(seg_14_11_local_g2_0_57897)
  );
  CascadeMux t20 (
    .I(net_16695),
    .O(net_16695_cascademuxed)
  );
  CascadeMux t200 (
    .I(net_44972),
    .O(net_44972_cascademuxed)
  );
  Span4Mux_h4 t2000 (
    .I(seg_12_11_sp4_v_t_42_46624),
    .O(seg_14_11_sp4_h_r_24_50314)
  );
  LocalMux t2001 (
    .I(seg_14_15_sp4_h_r_35_50809),
    .O(seg_14_15_local_g2_3_58392)
  );
  Span4Mux_h4 t2002 (
    .I(seg_12_15_sp4_v_t_46_47120),
    .O(seg_14_15_sp4_h_r_35_50809)
  );
  LocalMux t2003 (
    .I(seg_15_11_sp4_h_r_37_50314),
    .O(seg_15_11_local_g3_5_61740)
  );
  Span4Mux_h4 t2004 (
    .I(seg_12_11_sp4_v_t_42_46624),
    .O(seg_15_11_sp4_h_r_37_50314)
  );
  LocalMux t2005 (
    .I(seg_10_12_sp4_r_v_b_27_42666),
    .O(seg_10_12_local_g1_3_42692)
  );
  Span4Mux_v4 t2006 (
    .I(seg_11_14_sp4_v_t_42_43162),
    .O(seg_10_12_sp4_r_v_b_27_42666)
  );
  LocalMux t2007 (
    .I(seg_10_14_sp4_r_v_b_3_42666),
    .O(seg_10_14_local_g1_3_42938)
  );
  Span4Mux_v4 t2008 (
    .I(seg_11_14_sp4_v_t_42_43162),
    .O(seg_10_14_sp4_r_v_b_3_42666)
  );
  LocalMux t2009 (
    .I(seg_11_18_lutff_3_out_43381),
    .O(seg_11_18_local_g2_3_47269)
  );
  CascadeMux t201 (
    .I(net_45932),
    .O(net_45932_cascademuxed)
  );
  LocalMux t2010 (
    .I(seg_12_18_neigh_op_lft_4_43382),
    .O(seg_12_18_local_g0_4_51085)
  );
  LocalMux t2011 (
    .I(seg_11_18_lutff_5_out_43383),
    .O(seg_11_18_local_g2_5_47271)
  );
  LocalMux t2012 (
    .I(seg_15_18_sp4_h_r_2_62670),
    .O(seg_15_18_local_g1_2_62582)
  );
  Span4Mux_h4 t2013 (
    .I(seg_15_18_sp4_h_l_39_47348),
    .O(seg_15_18_sp4_h_r_2_62670)
  );
  LocalMux t2014 (
    .I(seg_14_18_sp4_h_r_41_47350),
    .O(seg_14_18_local_g2_1_58759)
  );
  LocalMux t2015 (
    .I(seg_12_19_neigh_op_lft_2_43503),
    .O(seg_12_19_local_g1_2_51214)
  );
  LocalMux t2016 (
    .I(seg_11_19_lutff_6_out_43507),
    .O(seg_11_19_local_g3_6_47403)
  );
  LocalMux t2017 (
    .I(seg_14_19_sp4_h_r_43_47475),
    .O(seg_14_19_local_g2_3_58884)
  );
  LocalMux t2018 (
    .I(seg_11_19_neigh_op_top_1_43625),
    .O(seg_11_19_local_g1_1_47382)
  );
  LocalMux t2019 (
    .I(seg_13_20_sp4_h_r_36_43760),
    .O(seg_13_20_local_g3_4_55186)
  );
  CascadeMux t202 (
    .I(net_45974),
    .O(net_45974_cascademuxed)
  );
  LocalMux t2020 (
    .I(seg_13_20_sp4_h_r_28_47596),
    .O(seg_13_20_local_g2_4_55178)
  );
  LocalMux t2021 (
    .I(seg_12_21_sp4_v_b_37_47726),
    .O(seg_12_21_local_g2_5_51471)
  );
  LocalMux t2022 (
    .I(seg_13_22_sp4_h_r_26_47840),
    .O(seg_13_22_local_g2_2_55422)
  );
  Span4Mux_h4 t2023 (
    .I(seg_11_22_sp4_v_t_44_44148),
    .O(seg_13_22_sp4_h_r_26_47840)
  );
  LocalMux t2024 (
    .I(seg_11_23_sp4_v_b_34_44028),
    .O(seg_11_23_local_g2_2_47883)
  );
  Span4Mux_v4 t2025 (
    .I(seg_11_25_sp4_v_t_47_44520),
    .O(seg_11_23_sp4_v_b_34_44028)
  );
  LocalMux t2026 (
    .I(seg_13_31_span4_horz_r_11_48881),
    .O(seg_13_31_local_g1_3_56535)
  );
  IoSpan4Mux t2027 (
    .I(seg_15_31_span4_vert_43_64169),
    .O(seg_13_31_span4_horz_r_11_48881)
  );
  Span4Mux_v4 t2028 (
    .I(seg_15_30_sp4_h_l_43_48824),
    .O(seg_15_31_span4_vert_43_64169)
  );
  LocalMux t2029 (
    .I(seg_11_8_neigh_op_rgt_1_45980),
    .O(seg_11_8_local_g2_1_46037)
  );
  CascadeMux t203 (
    .I(net_46061),
    .O(net_46061_cascademuxed)
  );
  LocalMux t2030 (
    .I(seg_12_8_lutff_1_out_45980),
    .O(seg_12_8_local_g3_1_49876)
  );
  LocalMux t2031 (
    .I(seg_11_9_neigh_op_bnr_5_45984),
    .O(seg_11_9_local_g0_5_46148)
  );
  LocalMux t2032 (
    .I(seg_12_8_lutff_5_out_45984),
    .O(seg_12_8_local_g2_5_49872)
  );
  LocalMux t2033 (
    .I(seg_9_8_sp4_h_r_15_34625),
    .O(seg_9_8_local_g1_7_38373)
  );
  Span4Mux_h4 t2034 (
    .I(seg_12_8_sp4_h_r_2_49949),
    .O(seg_9_8_sp4_h_r_15_34625)
  );
  LocalMux t2035 (
    .I(seg_12_8_sp4_r_v_b_3_49590),
    .O(seg_12_8_local_g1_3_49862)
  );
  Span4Mux_v4 t2036 (
    .I(seg_13_8_sp4_h_l_44_38463),
    .O(seg_12_8_sp4_r_v_b_3_49590)
  );
  LocalMux t2037 (
    .I(seg_12_11_lutff_0_out_46348),
    .O(seg_12_11_local_g0_0_50220)
  );
  LocalMux t2038 (
    .I(seg_12_12_neigh_op_bot_2_46350),
    .O(seg_12_12_local_g0_2_50345)
  );
  LocalMux t2039 (
    .I(seg_12_12_neigh_op_bot_5_46353),
    .O(seg_12_12_local_g0_5_50348)
  );
  CascadeMux t204 (
    .I(net_46067),
    .O(net_46067_cascademuxed)
  );
  LocalMux t2040 (
    .I(seg_12_11_lutff_6_out_46354),
    .O(seg_12_11_local_g0_6_50226)
  );
  LocalMux t2041 (
    .I(seg_14_11_sp4_h_r_26_50318),
    .O(seg_14_11_local_g2_2_57899)
  );
  LocalMux t2042 (
    .I(seg_16_12_sp4_h_r_47_54270),
    .O(seg_16_12_local_g2_7_65688)
  );
  Span4Mux_h4 t2043 (
    .I(seg_13_12_sp4_v_b_10_50091),
    .O(seg_16_12_sp4_h_r_47_54270)
  );
  LocalMux t2044 (
    .I(seg_11_12_neigh_op_rgt_1_46472),
    .O(seg_11_12_local_g2_1_46529)
  );
  LocalMux t2045 (
    .I(seg_13_12_neigh_op_lft_3_46474),
    .O(seg_13_12_local_g0_3_54177)
  );
  LocalMux t2046 (
    .I(seg_13_12_neigh_op_lft_4_46475),
    .O(seg_13_12_local_g1_4_54186)
  );
  LocalMux t2047 (
    .I(seg_11_12_neigh_op_rgt_5_46476),
    .O(seg_11_12_local_g2_5_46533)
  );
  LocalMux t2048 (
    .I(seg_13_12_neigh_op_lft_6_46477),
    .O(seg_13_12_local_g1_6_54188)
  );
  LocalMux t2049 (
    .I(seg_11_12_neigh_op_rgt_7_46478),
    .O(seg_11_12_local_g2_7_46535)
  );
  CascadeMux t205 (
    .I(net_46073),
    .O(net_46073_cascademuxed)
  );
  LocalMux t2050 (
    .I(seg_14_12_sp4_h_r_28_50443),
    .O(seg_14_12_local_g2_4_58024)
  );
  LocalMux t2051 (
    .I(seg_13_13_neigh_op_lft_0_46594),
    .O(seg_13_13_local_g1_0_54305)
  );
  LocalMux t2052 (
    .I(seg_11_13_neigh_op_rgt_1_46595),
    .O(seg_11_13_local_g2_1_46652)
  );
  LocalMux t2053 (
    .I(seg_11_13_neigh_op_rgt_2_46596),
    .O(seg_11_13_local_g2_2_46653)
  );
  LocalMux t2054 (
    .I(seg_13_13_neigh_op_lft_3_46597),
    .O(seg_13_13_local_g1_3_54308)
  );
  LocalMux t2055 (
    .I(seg_11_13_neigh_op_rgt_4_46598),
    .O(seg_11_13_local_g3_4_46663)
  );
  LocalMux t2056 (
    .I(seg_11_13_neigh_op_rgt_5_46599),
    .O(seg_11_13_local_g2_5_46656)
  );
  LocalMux t2057 (
    .I(seg_11_13_neigh_op_rgt_6_46600),
    .O(seg_11_13_local_g3_6_46665)
  );
  LocalMux t2058 (
    .I(seg_11_13_neigh_op_rgt_7_46601),
    .O(seg_11_13_local_g2_7_46658)
  );
  LocalMux t2059 (
    .I(seg_12_14_lutff_0_out_46717),
    .O(seg_12_14_local_g1_0_50597)
  );
  CascadeMux t206 (
    .I(net_46079),
    .O(net_46079_cascademuxed)
  );
  LocalMux t2060 (
    .I(seg_12_13_neigh_op_top_1_46718),
    .O(seg_12_13_local_g1_1_50475)
  );
  LocalMux t2061 (
    .I(seg_12_13_neigh_op_top_3_46720),
    .O(seg_12_13_local_g1_3_50477)
  );
  LocalMux t2062 (
    .I(seg_12_14_lutff_4_out_46721),
    .O(seg_12_14_local_g0_4_50593)
  );
  LocalMux t2063 (
    .I(seg_12_13_neigh_op_top_5_46722),
    .O(seg_12_13_local_g1_5_50479)
  );
  LocalMux t2064 (
    .I(seg_15_14_sp4_h_r_6_62182),
    .O(seg_15_14_local_g1_6_62094)
  );
  Span4Mux_h4 t2065 (
    .I(seg_15_14_sp4_h_l_38_46857),
    .O(seg_15_14_sp4_h_r_6_62182)
  );
  LocalMux t2066 (
    .I(seg_15_14_sp4_h_r_41_50689),
    .O(seg_15_14_local_g3_1_62105)
  );
  LocalMux t2067 (
    .I(seg_12_12_sp4_v_b_32_46504),
    .O(seg_12_12_local_g2_0_50359)
  );
  LocalMux t2068 (
    .I(seg_11_15_neigh_op_rgt_0_46840),
    .O(seg_11_15_local_g3_0_46905)
  );
  LocalMux t2069 (
    .I(seg_12_15_lutff_0_out_46840),
    .O(seg_12_15_local_g2_0_50728)
  );
  CascadeMux t207 (
    .I(net_46085),
    .O(net_46085_cascademuxed)
  );
  LocalMux t2070 (
    .I(seg_13_15_neigh_op_lft_4_46844),
    .O(seg_13_15_local_g1_4_54555)
  );
  LocalMux t2071 (
    .I(seg_13_15_neigh_op_lft_5_46845),
    .O(seg_13_15_local_g0_5_54548)
  );
  LocalMux t2072 (
    .I(seg_12_15_lutff_7_out_46847),
    .O(seg_12_15_local_g2_7_50735)
  );
  LocalMux t2073 (
    .I(seg_10_15_sp4_h_r_6_43152),
    .O(seg_10_15_local_g0_6_43056)
  );
  LocalMux t2074 (
    .I(seg_15_15_sp4_h_r_41_50812),
    .O(seg_15_15_local_g2_1_62220)
  );
  LocalMux t2075 (
    .I(seg_12_13_sp4_r_v_b_27_50451),
    .O(seg_12_13_local_g0_3_50469)
  );
  LocalMux t2076 (
    .I(seg_12_12_sp4_v_b_43_46625),
    .O(seg_12_12_local_g3_3_50370)
  );
  LocalMux t2077 (
    .I(seg_13_17_neigh_op_bnl_1_46964),
    .O(seg_13_17_local_g2_1_54806)
  );
  LocalMux t2078 (
    .I(seg_12_16_lutff_2_out_46965),
    .O(seg_12_16_local_g3_2_50861)
  );
  LocalMux t2079 (
    .I(seg_12_17_neigh_op_bot_4_46967),
    .O(seg_12_17_local_g0_4_50962)
  );
  CascadeMux t208 (
    .I(net_46091),
    .O(net_46091_cascademuxed)
  );
  LocalMux t2080 (
    .I(seg_13_15_neigh_op_tnl_5_46968),
    .O(seg_13_15_local_g3_5_54572)
  );
  LocalMux t2081 (
    .I(seg_13_15_neigh_op_tnl_6_46969),
    .O(seg_13_15_local_g2_6_54565)
  );
  LocalMux t2082 (
    .I(seg_14_16_sp4_h_r_32_50939),
    .O(seg_14_16_local_g3_0_58520)
  );
  LocalMux t2083 (
    .I(seg_13_17_neigh_op_lft_0_47086),
    .O(seg_13_17_local_g1_0_54797)
  );
  LocalMux t2084 (
    .I(seg_12_16_neigh_op_top_1_47087),
    .O(seg_12_16_local_g0_1_50836)
  );
  LocalMux t2085 (
    .I(seg_12_17_lutff_1_out_47087),
    .O(seg_12_17_local_g1_1_50967)
  );
  LocalMux t2086 (
    .I(seg_13_17_neigh_op_lft_3_47089),
    .O(seg_13_17_local_g0_3_54792)
  );
  LocalMux t2087 (
    .I(seg_12_17_lutff_5_out_47091),
    .O(seg_12_17_local_g1_5_50971)
  );
  LocalMux t2088 (
    .I(seg_13_17_neigh_op_lft_6_47092),
    .O(seg_13_17_local_g0_6_54795)
  );
  LocalMux t2089 (
    .I(seg_16_15_sp4_v_b_28_62191),
    .O(seg_16_15_local_g3_4_66062)
  );
  CascadeMux t209 (
    .I(net_46097),
    .O(net_46097_cascademuxed)
  );
  Span4Mux_v4 t2090 (
    .I(seg_16_17_sp4_h_l_47_51054),
    .O(seg_16_15_sp4_v_b_28_62191)
  );
  LocalMux t2091 (
    .I(seg_12_18_lutff_2_out_47211),
    .O(seg_12_18_local_g2_2_51099)
  );
  LocalMux t2092 (
    .I(seg_12_18_lutff_5_out_47214),
    .O(seg_12_18_local_g0_5_51086)
  );
  LocalMux t2093 (
    .I(seg_13_19_neigh_op_bnl_7_47216),
    .O(seg_13_19_local_g3_7_55066)
  );
  LocalMux t2094 (
    .I(seg_19_18_sp4_h_r_45_66507),
    .O(seg_19_18_local_g2_5_77558)
  );
  Span4Mux_h4 t2095 (
    .I(seg_16_18_sp4_h_l_37_51175),
    .O(seg_19_18_sp4_h_r_45_66507)
  );
  LocalMux t2096 (
    .I(seg_18_17_sp4_r_v_b_21_73811),
    .O(seg_18_17_local_g3_5_73971)
  );
  Span4Mux_v4 t2097 (
    .I(seg_19_18_sp4_h_l_45_62676),
    .O(seg_18_17_sp4_r_v_b_21_73811)
  );
  Span4Mux_h4 t2098 (
    .I(seg_15_18_sp4_h_l_40_47351),
    .O(seg_19_18_sp4_h_l_45_62676)
  );
  LocalMux t2099 (
    .I(seg_12_19_lutff_3_out_47335),
    .O(seg_12_19_local_g3_3_51231)
  );
  CascadeMux t21 (
    .I(net_17280),
    .O(net_17280_cascademuxed)
  );
  CascadeMux t210 (
    .I(net_46202),
    .O(net_46202_cascademuxed)
  );
  LocalMux t2100 (
    .I(seg_12_19_lutff_4_out_47336),
    .O(seg_12_19_local_g1_4_51216)
  );
  LocalMux t2101 (
    .I(seg_12_19_lutff_6_out_47338),
    .O(seg_12_19_local_g0_6_51210)
  );
  LocalMux t2102 (
    .I(seg_12_18_neigh_op_top_7_47339),
    .O(seg_12_18_local_g0_7_51088)
  );
  LocalMux t2103 (
    .I(seg_19_18_sp4_r_v_b_18_77425),
    .O(seg_19_18_local_g3_2_77563)
  );
  Span4Mux_v4 t2104 (
    .I(seg_20_19_sp4_h_l_42_66629),
    .O(seg_19_18_sp4_r_v_b_18_77425)
  );
  Span4Mux_h4 t2105 (
    .I(seg_16_19_sp4_h_l_41_51304),
    .O(seg_20_19_sp4_h_l_42_66629)
  );
  LocalMux t2106 (
    .I(seg_17_18_sp4_h_r_5_70335),
    .O(seg_17_18_local_g1_5_70247)
  );
  Span4Mux_h4 t2107 (
    .I(seg_17_18_sp4_h_l_40_55013),
    .O(seg_17_18_sp4_h_r_5_70335)
  );
  Span4Mux_h4 t2108 (
    .I(seg_13_18_sp4_v_t_37_51311),
    .O(seg_17_18_sp4_h_l_40_55013)
  );
  LocalMux t2109 (
    .I(seg_12_19_neigh_op_top_1_47456),
    .O(seg_12_19_local_g1_1_51213)
  );
  CascadeMux t211 (
    .I(net_46208),
    .O(net_46208_cascademuxed)
  );
  LocalMux t2110 (
    .I(seg_12_21_lutff_2_out_47580),
    .O(seg_12_21_local_g1_2_51460)
  );
  LocalMux t2111 (
    .I(seg_13_20_neigh_op_tnl_2_47580),
    .O(seg_13_20_local_g2_2_55176)
  );
  LocalMux t2112 (
    .I(seg_12_21_lutff_6_out_47584),
    .O(seg_12_21_local_g0_6_51456)
  );
  LocalMux t2113 (
    .I(seg_14_11_sp12_h_r_4_50310),
    .O(seg_14_11_local_g0_4_57885)
  );
  Span12Mux_h12 t2114 (
    .I(seg_12_11_sp12_v_t_23_50313),
    .O(seg_14_11_sp12_h_r_4_50310)
  );
  LocalMux t2115 (
    .I(seg_16_20_sp4_v_b_19_62685),
    .O(seg_16_20_local_g1_3_66660)
  );
  Span4Mux_v4 t2116 (
    .I(seg_16_21_sp4_h_l_37_51544),
    .O(seg_16_20_sp4_v_b_19_62685)
  );
  LocalMux t2117 (
    .I(seg_12_21_sp4_h_r_19_47721),
    .O(seg_12_21_local_g1_3_51461)
  );
  Span4Mux_h4 t2118 (
    .I(seg_15_21_sp4_h_r_3_63040),
    .O(seg_12_21_sp4_h_r_19_47721)
  );
  Span4Mux_h4 t2119 (
    .I(seg_15_21_sp4_h_l_38_47718),
    .O(seg_15_21_sp4_h_r_3_63040)
  );
  CascadeMux t212 (
    .I(net_46214),
    .O(net_46214_cascademuxed)
  );
  LocalMux t2120 (
    .I(seg_11_19_sp4_v_b_34_43536),
    .O(seg_11_19_local_g2_2_47391)
  );
  Span4Mux_v4 t2121 (
    .I(seg_11_21_sp4_h_r_5_47720),
    .O(seg_11_19_sp4_v_b_34_43536)
  );
  LocalMux t2122 (
    .I(seg_14_12_sp4_r_v_b_14_57866),
    .O(seg_14_12_local_g2_6_58026)
  );
  Span4Mux_v4 t2123 (
    .I(seg_15_13_sp4_v_t_37_58357),
    .O(seg_14_12_sp4_r_v_b_14_57866)
  );
  Span4Mux_v4 t2124 (
    .I(seg_15_17_sp4_v_t_44_58856),
    .O(seg_15_13_sp4_v_t_37_58357)
  );
  Span4Mux_v4 t2125 (
    .I(seg_15_21_sp4_h_l_44_47724),
    .O(seg_15_17_sp4_v_t_44_58856)
  );
  LocalMux t2126 (
    .I(seg_14_15_sp4_r_v_b_29_58360),
    .O(seg_14_15_local_g1_5_58386)
  );
  Span4Mux_v4 t2127 (
    .I(seg_15_17_sp4_v_t_44_58856),
    .O(seg_14_15_sp4_r_v_b_29_58360)
  );
  LocalMux t2128 (
    .I(seg_14_16_sp4_r_v_b_13_58357),
    .O(seg_14_16_local_g2_5_58517)
  );
  Span4Mux_v4 t2129 (
    .I(seg_15_17_sp4_v_t_44_58856),
    .O(seg_14_16_sp4_r_v_b_13_58357)
  );
  CascadeMux t213 (
    .I(net_46220),
    .O(net_46220_cascademuxed)
  );
  LocalMux t2130 (
    .I(seg_14_19_sp4_r_v_b_33_58856),
    .O(seg_14_19_local_g0_2_58867)
  );
  Span4Mux_v4 t2131 (
    .I(seg_15_21_sp4_h_l_44_47724),
    .O(seg_14_19_sp4_r_v_b_33_58856)
  );
  LocalMux t2132 (
    .I(seg_14_20_sp4_r_v_b_20_58856),
    .O(seg_14_20_local_g3_4_59016)
  );
  Span4Mux_v4 t2133 (
    .I(seg_15_21_sp4_h_l_44_47724),
    .O(seg_14_20_sp4_r_v_b_20_58856)
  );
  LocalMux t2134 (
    .I(seg_15_10_sp4_v_b_38_57866),
    .O(seg_15_10_local_g2_6_61610)
  );
  Span4Mux_v4 t2135 (
    .I(seg_15_13_sp4_v_t_37_58357),
    .O(seg_15_10_sp4_v_b_38_57866)
  );
  LocalMux t2136 (
    .I(seg_15_16_sp4_v_b_16_58360),
    .O(seg_15_16_local_g1_0_62334)
  );
  Span4Mux_v4 t2137 (
    .I(seg_15_17_sp4_v_t_44_58856),
    .O(seg_15_16_sp4_v_b_16_58360)
  );
  LocalMux t2138 (
    .I(seg_15_19_sp4_v_b_33_58856),
    .O(seg_15_19_local_g3_1_62720)
  );
  Span4Mux_v4 t2139 (
    .I(seg_15_21_sp4_h_l_44_47724),
    .O(seg_15_19_sp4_v_b_33_58856)
  );
  CascadeMux t214 (
    .I(net_46301),
    .O(net_46301_cascademuxed)
  );
  LocalMux t2140 (
    .I(seg_14_12_sp4_v_b_18_54040),
    .O(seg_14_12_local_g0_2_58006)
  );
  Span4Mux_v4 t2141 (
    .I(seg_14_13_sp4_v_t_41_54531),
    .O(seg_14_12_sp4_v_b_18_54040)
  );
  Span4Mux_v4 t2142 (
    .I(seg_14_17_sp4_v_t_45_55027),
    .O(seg_14_13_sp4_v_t_41_54531)
  );
  Span4Mux_v4 t2143 (
    .I(seg_14_21_sp4_h_l_45_43892),
    .O(seg_14_17_sp4_v_t_45_55027)
  );
  LocalMux t2144 (
    .I(seg_16_19_sp4_v_b_28_62683),
    .O(seg_16_19_local_g2_4_66546)
  );
  Span4Mux_v4 t2145 (
    .I(seg_16_21_sp4_h_l_41_51550),
    .O(seg_16_19_sp4_v_b_28_62683)
  );
  LocalMux t2146 (
    .I(seg_16_20_sp4_v_b_17_62683),
    .O(seg_16_20_local_g0_1_66650)
  );
  Span4Mux_v4 t2147 (
    .I(seg_16_21_sp4_h_l_41_51550),
    .O(seg_16_20_sp4_v_b_17_62683)
  );
  LocalMux t2148 (
    .I(seg_13_12_sp4_v_b_18_50209),
    .O(seg_13_12_local_g0_2_54176)
  );
  Span4Mux_v4 t2149 (
    .I(seg_13_13_sp4_v_t_41_50700),
    .O(seg_13_12_sp4_v_b_18_50209)
  );
  CascadeMux t215 (
    .I(net_46319),
    .O(net_46319_cascademuxed)
  );
  Span4Mux_v4 t2150 (
    .I(seg_13_17_sp4_v_t_36_51187),
    .O(seg_13_13_sp4_v_t_41_50700)
  );
  LocalMux t2151 (
    .I(seg_13_20_sp4_v_b_19_51194),
    .O(seg_13_20_local_g1_3_55169)
  );
  Span4Mux_v4 t2152 (
    .I(seg_13_21_sp4_h_r_1_55376),
    .O(seg_13_20_sp4_v_b_19_51194)
  );
  Span4Mux_h4 t2153 (
    .I(seg_13_21_sp4_v_b_1_51187),
    .O(seg_13_21_sp4_h_r_1_55376)
  );
  LocalMux t2154 (
    .I(seg_11_14_sp4_h_r_34_39192),
    .O(seg_11_14_local_g2_2_46776)
  );
  Span4Mux_h4 t2155 (
    .I(seg_13_14_sp4_v_t_41_50823),
    .O(seg_11_14_sp4_h_r_34_39192)
  );
  Span4Mux_v4 t2156 (
    .I(seg_13_18_sp4_v_t_41_51315),
    .O(seg_13_14_sp4_v_t_41_50823)
  );
  LocalMux t2157 (
    .I(seg_11_18_sp4_h_r_34_39684),
    .O(seg_11_18_local_g2_2_47268)
  );
  Span4Mux_h4 t2158 (
    .I(seg_13_18_sp4_v_t_41_51315),
    .O(seg_11_18_sp4_h_r_34_39684)
  );
  LocalMux t2159 (
    .I(seg_13_11_sp4_v_b_42_50332),
    .O(seg_13_11_local_g2_2_54069)
  );
  CascadeMux t216 (
    .I(net_46331),
    .O(net_46331_cascademuxed)
  );
  Span4Mux_v4 t2160 (
    .I(seg_13_14_sp4_v_t_42_50824),
    .O(seg_13_11_sp4_v_b_42_50332)
  );
  Span4Mux_v4 t2161 (
    .I(seg_13_18_sp4_v_t_41_51315),
    .O(seg_13_14_sp4_v_t_42_50824)
  );
  LocalMux t2162 (
    .I(seg_14_10_sp4_h_r_22_54025),
    .O(seg_14_10_local_g0_6_57764)
  );
  Span4Mux_h4 t2163 (
    .I(seg_13_10_sp4_v_t_46_50336),
    .O(seg_14_10_sp4_h_r_22_54025)
  );
  Span4Mux_v4 t2164 (
    .I(seg_13_14_sp4_v_t_45_50827),
    .O(seg_13_10_sp4_v_t_46_50336)
  );
  Span4Mux_v4 t2165 (
    .I(seg_13_18_sp4_v_t_45_51319),
    .O(seg_13_14_sp4_v_t_45_50827)
  );
  LocalMux t2166 (
    .I(seg_15_18_sp4_h_r_25_55007),
    .O(seg_15_18_local_g2_1_62589)
  );
  Span4Mux_h4 t2167 (
    .I(seg_13_18_sp4_v_t_45_51319),
    .O(seg_15_18_sp4_h_r_25_55007)
  );
  LocalMux t2168 (
    .I(seg_12_11_sp4_r_v_b_32_50212),
    .O(seg_12_11_local_g0_3_50223)
  );
  Span4Mux_v4 t2169 (
    .I(seg_13_13_sp4_v_t_40_50699),
    .O(seg_12_11_sp4_r_v_b_32_50212)
  );
  CascadeMux t217 (
    .I(net_46337),
    .O(net_46337_cascademuxed)
  );
  Span4Mux_v4 t2170 (
    .I(seg_13_17_sp4_v_t_40_51191),
    .O(seg_13_13_sp4_v_t_40_50699)
  );
  LocalMux t2171 (
    .I(seg_12_14_sp4_r_v_b_40_50699),
    .O(seg_12_14_local_g3_0_50613)
  );
  Span4Mux_v4 t2172 (
    .I(seg_13_17_sp4_v_t_40_51191),
    .O(seg_12_14_sp4_r_v_b_40_50699)
  );
  LocalMux t2173 (
    .I(seg_13_12_sp4_v_b_21_50212),
    .O(seg_13_12_local_g1_5_54187)
  );
  Span4Mux_v4 t2174 (
    .I(seg_13_13_sp4_v_t_40_50699),
    .O(seg_13_12_sp4_v_b_21_50212)
  );
  LocalMux t2175 (
    .I(seg_13_13_sp4_h_r_5_54398),
    .O(seg_13_13_local_g0_5_54302)
  );
  Span4Mux_h4 t2176 (
    .I(seg_13_13_sp4_v_t_40_50699),
    .O(seg_13_13_sp4_h_r_5_54398)
  );
  LocalMux t2177 (
    .I(seg_13_14_sp4_v_b_40_50699),
    .O(seg_13_14_local_g3_0_54444)
  );
  Span4Mux_v4 t2178 (
    .I(seg_13_17_sp4_v_t_40_51191),
    .O(seg_13_14_sp4_v_b_40_50699)
  );
  LocalMux t2179 (
    .I(seg_13_19_sp4_v_b_29_51191),
    .O(seg_13_19_local_g2_5_55056)
  );
  CascadeMux t218 (
    .I(net_46436),
    .O(net_46436_cascademuxed)
  );
  LocalMux t2180 (
    .I(seg_14_13_sp4_h_r_16_54398),
    .O(seg_14_13_local_g1_0_58135)
  );
  Span4Mux_h4 t2181 (
    .I(seg_13_13_sp4_v_t_40_50699),
    .O(seg_14_13_sp4_h_r_16_54398)
  );
  LocalMux t2182 (
    .I(seg_15_17_sp4_h_r_29_54890),
    .O(seg_15_17_local_g2_5_62470)
  );
  Span4Mux_h4 t2183 (
    .I(seg_13_17_sp4_v_t_40_51191),
    .O(seg_15_17_sp4_h_r_29_54890)
  );
  LocalMux t2184 (
    .I(seg_16_12_sp4_r_v_b_16_65529),
    .O(seg_16_12_local_g3_0_65689)
  );
  Span4Mux_v4 t2185 (
    .I(seg_17_13_sp4_h_l_40_54398),
    .O(seg_16_12_sp4_r_v_b_16_65529)
  );
  Span4Mux_h4 t2186 (
    .I(seg_13_13_sp4_v_t_40_50699),
    .O(seg_17_13_sp4_h_l_40_54398)
  );
  LocalMux t2187 (
    .I(seg_16_16_sp4_r_v_b_16_66021),
    .O(seg_16_16_local_g3_0_66181)
  );
  Span4Mux_v4 t2188 (
    .I(seg_17_17_sp4_h_l_40_54890),
    .O(seg_16_16_sp4_r_v_b_16_66021)
  );
  Span4Mux_h4 t2189 (
    .I(seg_13_17_sp4_v_t_40_51191),
    .O(seg_17_17_sp4_h_l_40_54890)
  );
  LocalMux t2190 (
    .I(seg_12_13_sp4_h_r_43_39075),
    .O(seg_12_13_local_g3_3_50493)
  );
  Span4Mux_h4 t2191 (
    .I(seg_13_13_sp4_v_t_37_50696),
    .O(seg_12_13_sp4_h_r_43_39075)
  );
  Span4Mux_v4 t2192 (
    .I(seg_13_17_sp4_v_t_44_51195),
    .O(seg_13_13_sp4_v_t_37_50696)
  );
  LocalMux t2193 (
    .I(seg_11_15_sp4_r_v_b_27_46866),
    .O(seg_11_15_local_g1_3_46892)
  );
  Span4Mux_v4 t2194 (
    .I(seg_12_17_sp4_v_t_37_47357),
    .O(seg_11_15_sp4_r_v_b_27_46866)
  );
  LocalMux t2195 (
    .I(seg_12_11_sp4_v_b_35_46382),
    .O(seg_12_11_local_g3_3_50247)
  );
  Span4Mux_v4 t2196 (
    .I(seg_12_13_sp4_v_t_38_46866),
    .O(seg_12_11_sp4_v_b_35_46382)
  );
  Span4Mux_v4 t2197 (
    .I(seg_12_17_sp4_v_t_37_47357),
    .O(seg_12_13_sp4_v_t_38_46866)
  );
  LocalMux t2198 (
    .I(seg_14_13_sp4_h_r_27_50565),
    .O(seg_14_13_local_g3_3_58154)
  );
  Span4Mux_h4 t2199 (
    .I(seg_12_13_sp4_v_t_38_46866),
    .O(seg_14_13_sp4_h_r_27_50565)
  );
  CascadeMux t22 (
    .I(net_17286),
    .O(net_17286_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t220 (
    .carryinitin(),
    .carryinitout(t219)
  );
  LocalMux t2200 (
    .I(seg_13_14_sp4_h_r_19_50691),
    .O(seg_13_14_local_g1_3_54431)
  );
  Span4Mux_h4 t2201 (
    .I(seg_12_14_sp4_v_t_36_46987),
    .O(seg_13_14_sp4_h_r_19_50691)
  );
  Span4Mux_v4 t2202 (
    .I(seg_12_18_sp4_v_t_40_47483),
    .O(seg_12_14_sp4_v_t_36_46987)
  );
  LocalMux t2203 (
    .I(seg_11_12_sp4_r_v_b_14_46374),
    .O(seg_11_12_local_g2_6_46534)
  );
  Span4Mux_v4 t2204 (
    .I(seg_12_13_sp4_v_t_42_46870),
    .O(seg_11_12_sp4_r_v_b_14_46374)
  );
  Span4Mux_v4 t2205 (
    .I(seg_12_17_sp4_v_t_41_47361),
    .O(seg_12_13_sp4_v_t_42_46870)
  );
  LocalMux t2206 (
    .I(seg_11_13_sp4_r_v_b_3_46374),
    .O(seg_11_13_local_g1_3_46646)
  );
  Span4Mux_v4 t2207 (
    .I(seg_12_13_sp4_v_t_42_46870),
    .O(seg_11_13_sp4_r_v_b_3_46374)
  );
  LocalMux t2208 (
    .I(seg_11_14_sp4_r_v_b_42_46870),
    .O(seg_11_14_local_g3_2_46784)
  );
  Span4Mux_v4 t2209 (
    .I(seg_12_17_sp4_v_t_41_47361),
    .O(seg_11_14_sp4_r_v_b_42_46870)
  );
  CascadeMux t221 (
    .I(net_46553),
    .O(net_46553_cascademuxed)
  );
  LocalMux t2210 (
    .I(seg_11_18_sp4_r_v_b_41_47361),
    .O(seg_11_18_local_g3_1_47275)
  );
  LocalMux t2211 (
    .I(seg_11_19_sp4_r_v_b_28_47361),
    .O(seg_11_19_local_g0_4_47377)
  );
  LocalMux t2212 (
    .I(seg_12_11_sp4_v_b_27_46374),
    .O(seg_12_11_local_g2_3_50239)
  );
  Span4Mux_v4 t2213 (
    .I(seg_12_13_sp4_v_t_42_46870),
    .O(seg_12_11_sp4_v_b_27_46374)
  );
  LocalMux t2214 (
    .I(seg_12_14_sp4_v_b_42_46870),
    .O(seg_12_14_local_g3_2_50615)
  );
  Span4Mux_v4 t2215 (
    .I(seg_12_17_sp4_v_t_41_47361),
    .O(seg_12_14_sp4_v_b_42_46870)
  );
  LocalMux t2216 (
    .I(seg_12_15_sp4_v_b_31_46870),
    .O(seg_12_15_local_g3_7_50743)
  );
  Span4Mux_v4 t2217 (
    .I(seg_12_17_sp4_v_t_41_47361),
    .O(seg_12_15_sp4_v_b_31_46870)
  );
  LocalMux t2218 (
    .I(seg_12_18_sp4_v_b_41_47361),
    .O(seg_12_18_local_g3_1_51106)
  );
  LocalMux t2219 (
    .I(seg_12_12_sp4_v_b_19_46379),
    .O(seg_12_12_local_g1_3_50354)
  );
  CascadeMux t222 (
    .I(net_46565),
    .O(net_46565_cascademuxed)
  );
  Span4Mux_v4 t2220 (
    .I(seg_12_13_sp4_h_r_1_50561),
    .O(seg_12_12_sp4_v_b_19_46379)
  );
  Span4Mux_h4 t2221 (
    .I(seg_12_13_sp4_v_t_45_46873),
    .O(seg_12_13_sp4_h_r_1_50561)
  );
  Span4Mux_v4 t2222 (
    .I(seg_12_17_sp4_v_t_45_47365),
    .O(seg_12_13_sp4_v_t_45_46873)
  );
  LocalMux t2223 (
    .I(seg_12_14_sp4_v_b_43_46871),
    .O(seg_12_14_local_g3_3_50616)
  );
  Span4Mux_v4 t2224 (
    .I(seg_12_17_sp4_h_r_1_51053),
    .O(seg_12_14_sp4_v_b_43_46871)
  );
  Span4Mux_h4 t2225 (
    .I(seg_12_17_sp4_v_t_45_47365),
    .O(seg_12_17_sp4_h_r_1_51053)
  );
  LocalMux t2226 (
    .I(seg_14_2_sp4_v_b_14_52911),
    .O(seg_14_2_local_g0_6_56780)
  );
  Span4Mux_v4 t2227 (
    .I(seg_14_3_sp4_v_t_42_53302),
    .O(seg_14_2_sp4_v_b_14_52911)
  );
  Span4Mux_v4 t2228 (
    .I(seg_14_7_sp4_v_t_41_53793),
    .O(seg_14_3_sp4_v_t_42_53302)
  );
  Span4Mux_v4 t2229 (
    .I(seg_14_11_sp4_v_t_45_54289),
    .O(seg_14_7_sp4_v_t_41_53793)
  );
  CascadeMux t223 (
    .I(net_46571),
    .O(net_46571_cascademuxed)
  );
  Span4Mux_v4 t2230 (
    .I(seg_14_15_sp4_v_t_40_54776),
    .O(seg_14_11_sp4_v_t_45_54289)
  );
  Span4Mux_v4 t2231 (
    .I(seg_14_19_sp4_v_t_39_55267),
    .O(seg_14_15_sp4_v_t_40_54776)
  );
  Span4Mux_v4 t2232 (
    .I(seg_14_23_sp4_h_l_45_44138),
    .O(seg_14_19_sp4_v_t_39_55267)
  );
  LocalMux t2233 (
    .I(seg_14_4_sp4_v_b_42_53302),
    .O(seg_14_4_local_g3_2_57046)
  );
  Span4Mux_v4 t2234 (
    .I(seg_14_7_sp4_v_t_41_53793),
    .O(seg_14_4_sp4_v_b_42_53302)
  );
  LocalMux t2235 (
    .I(seg_13_3_sp4_h_r_11_53164),
    .O(seg_13_3_local_g1_3_53078)
  );
  Span4Mux_h4 t2236 (
    .I(seg_13_3_sp4_v_t_46_49475),
    .O(seg_13_3_sp4_h_r_11_53164)
  );
  Span4Mux_v4 t2237 (
    .I(seg_13_7_sp4_v_t_38_49959),
    .O(seg_13_3_sp4_v_t_46_49475)
  );
  Span4Mux_v4 t2238 (
    .I(seg_13_11_sp4_v_t_42_50455),
    .O(seg_13_7_sp4_v_t_38_49959)
  );
  Span4Mux_v4 t2239 (
    .I(seg_13_15_sp4_v_t_41_50946),
    .O(seg_13_11_sp4_v_t_42_50455)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t224 (
    .carryinitin(net_50417),
    .carryinitout(net_50461)
  );
  Span4Mux_v4 t2240 (
    .I(seg_13_19_sp4_v_t_36_51433),
    .O(seg_13_15_sp4_v_t_41_50946)
  );
  LocalMux t2241 (
    .I(seg_15_3_sp4_h_r_35_53164),
    .O(seg_15_3_local_g3_3_60754)
  );
  Span4Mux_h4 t2242 (
    .I(seg_13_3_sp4_v_t_46_49475),
    .O(seg_15_3_sp4_h_r_35_53164)
  );
  LocalMux t2243 (
    .I(seg_16_2_sp4_r_v_b_19_64406),
    .O(seg_16_2_local_g3_3_64462)
  );
  Span4Mux_v4 t2244 (
    .I(seg_17_3_sp4_h_l_43_53169),
    .O(seg_16_2_sp4_r_v_b_19_64406)
  );
  Span4Mux_h4 t2245 (
    .I(seg_13_3_sp4_v_t_43_49472),
    .O(seg_17_3_sp4_h_l_43_53169)
  );
  Span4Mux_v4 t2246 (
    .I(seg_13_7_sp4_v_t_38_49959),
    .O(seg_13_3_sp4_v_t_43_49472)
  );
  LocalMux t2247 (
    .I(seg_15_2_sp4_r_v_b_16_60573),
    .O(seg_15_2_local_g3_0_60628)
  );
  Span4Mux_v4 t2248 (
    .I(seg_16_3_sp4_h_l_46_49333),
    .O(seg_15_2_sp4_r_v_b_16_60573)
  );
  Span4Mux_h4 t2249 (
    .I(seg_12_3_sp4_v_t_43_45641),
    .O(seg_16_3_sp4_h_l_46_49333)
  );
  CascadeMux t225 (
    .I(net_46670),
    .O(net_46670_cascademuxed)
  );
  Span4Mux_v4 t2250 (
    .I(seg_12_7_sp4_v_t_43_46133),
    .O(seg_12_3_sp4_v_t_43_45641)
  );
  Span4Mux_v4 t2251 (
    .I(seg_12_11_sp4_v_t_38_46620),
    .O(seg_12_7_sp4_v_t_43_46133)
  );
  Span4Mux_v4 t2252 (
    .I(seg_12_15_sp4_v_t_38_47112),
    .O(seg_12_11_sp4_v_t_38_46620)
  );
  Span4Mux_v4 t2253 (
    .I(seg_12_19_sp4_v_t_37_47603),
    .O(seg_12_15_sp4_v_t_38_47112)
  );
  LocalMux t2254 (
    .I(seg_12_27_lutff_2_out_48318),
    .O(seg_12_27_local_g2_2_52206)
  );
  LocalMux t2255 (
    .I(seg_12_27_lutff_3_out_48319),
    .O(seg_12_27_local_g2_3_52207)
  );
  LocalMux t2256 (
    .I(seg_13_27_neigh_op_lft_4_48320),
    .O(seg_13_27_local_g1_4_56031)
  );
  LocalMux t2257 (
    .I(seg_13_27_neigh_op_lft_5_48321),
    .O(seg_13_27_local_g0_5_56024)
  );
  LocalMux t2258 (
    .I(seg_12_27_lutff_6_out_48322),
    .O(seg_12_27_local_g3_6_52218)
  );
  LocalMux t2259 (
    .I(seg_13_27_neigh_op_lft_6_48322),
    .O(seg_13_27_local_g0_6_56025)
  );
  CascadeMux t226 (
    .I(net_46676),
    .O(net_46676_cascademuxed)
  );
  LocalMux t2260 (
    .I(seg_12_27_lutff_7_out_48323),
    .O(seg_12_27_local_g0_7_52195)
  );
  LocalMux t2261 (
    .I(seg_13_27_neigh_op_lft_7_48323),
    .O(seg_13_27_local_g1_7_56034)
  );
  LocalMux t2262 (
    .I(seg_14_27_sp4_h_r_36_48452),
    .O(seg_14_27_local_g2_4_59869)
  );
  LocalMux t2263 (
    .I(seg_14_27_sp4_h_r_38_48456),
    .O(seg_14_27_local_g3_6_59879)
  );
  LocalMux t2264 (
    .I(seg_12_27_neigh_op_top_1_48440),
    .O(seg_12_27_local_g1_1_52197)
  );
  LocalMux t2265 (
    .I(seg_12_28_lutff_1_out_48440),
    .O(seg_12_28_local_g3_1_52336)
  );
  LocalMux t2266 (
    .I(seg_13_27_neigh_op_tnl_1_48440),
    .O(seg_13_27_local_g2_1_56036)
  );
  LocalMux t2267 (
    .I(seg_12_28_lutff_2_out_48441),
    .O(seg_12_28_local_g1_2_52321)
  );
  LocalMux t2268 (
    .I(seg_14_27_sp4_r_v_b_18_59715),
    .O(seg_14_27_local_g3_2_59875)
  );
  Span4Mux_v4 t2269 (
    .I(seg_15_28_sp4_h_l_42_48583),
    .O(seg_14_27_sp4_r_v_b_18_59715)
  );
  CascadeMux t227 (
    .I(net_46682),
    .O(net_46682_cascademuxed)
  );
  GlobalMux t2270 (
    .I(seg_13_0_local_g1_4_52735_i3),
    .O(seg_2_8_glb_netwk_0_5)
  );
  gio2CtrlBuf t2271 (
    .I(seg_13_0_local_g1_4_52735_i2),
    .O(seg_13_0_local_g1_4_52735_i3)
  );
  ICE_GB t2272 (
    .GLOBALBUFFEROUTPUT(seg_13_0_local_g1_4_52735_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_13_0_local_g1_4_52735_i1)
  );
  IoInMux t2273 (
    .I(seg_13_0_local_g1_4_52735),
    .O(seg_13_0_local_g1_4_52735_i1)
  );
  LocalMux t2274 (
    .I(seg_13_0_span4_horz_r_4_48940),
    .O(seg_13_0_local_g1_4_52735)
  );
  IoSpan4Mux t2275 (
    .I(seg_12_0_span4_vert_25_45247),
    .O(seg_13_0_span4_horz_r_4_48940)
  );
  Span4Mux_v4 t2276 (
    .I(seg_12_3_sp4_v_t_36_45634),
    .O(seg_12_0_span4_vert_25_45247)
  );
  Span4Mux_v4 t2277 (
    .I(seg_12_7_sp4_v_t_47_46137),
    .O(seg_12_3_sp4_v_t_36_45634)
  );
  Sp12to4 t2278 (
    .I(seg_12_10_sp12_v_b_23_50067),
    .O(seg_12_7_sp4_v_t_47_46137)
  );
  Span12Mux_v12 t2279 (
    .I(seg_12_21_sp12_v_t_23_51543),
    .O(seg_12_10_sp12_v_b_23_50067)
  );
  CascadeMux t228 (
    .I(net_46688),
    .O(net_46688_cascademuxed)
  );
  LocalMux t2280 (
    .I(seg_14_3_neigh_op_lft_7_49202),
    .O(seg_14_3_local_g1_7_56912)
  );
  LocalMux t2281 (
    .I(seg_14_3_sp4_v_b_19_52929),
    .O(seg_14_3_local_g1_3_56908)
  );
  LocalMux t2282 (
    .I(seg_14_4_neigh_op_lft_2_49320),
    .O(seg_14_4_local_g1_2_57030)
  );
  LocalMux t2283 (
    .I(seg_14_4_neigh_op_lft_3_49321),
    .O(seg_14_4_local_g0_3_57023)
  );
  LocalMux t2284 (
    .I(seg_13_4_lutff_4_out_49322),
    .O(seg_13_4_local_g0_4_53194)
  );
  LocalMux t2285 (
    .I(seg_13_4_lutff_5_out_49323),
    .O(seg_13_4_local_g2_5_53211)
  );
  LocalMux t2286 (
    .I(seg_13_3_neigh_op_top_6_49324),
    .O(seg_13_3_local_g0_6_53073)
  );
  LocalMux t2287 (
    .I(seg_13_4_lutff_6_out_49324),
    .O(seg_13_4_local_g1_6_53204)
  );
  LocalMux t2288 (
    .I(seg_13_3_neigh_op_top_7_49325),
    .O(seg_13_3_local_g0_7_53074)
  );
  LocalMux t2289 (
    .I(seg_13_4_lutff_7_out_49325),
    .O(seg_13_4_local_g2_7_53213)
  );
  CascadeMux t229 (
    .I(net_46694),
    .O(net_46694_cascademuxed)
  );
  LocalMux t2290 (
    .I(seg_13_9_neigh_op_bot_2_49812),
    .O(seg_13_9_local_g0_2_53807)
  );
  LocalMux t2291 (
    .I(seg_14_8_neigh_op_lft_3_49813),
    .O(seg_14_8_local_g0_3_57515)
  );
  LocalMux t2292 (
    .I(seg_13_9_neigh_op_bot_4_49814),
    .O(seg_13_9_local_g0_4_53809)
  );
  LocalMux t2293 (
    .I(seg_13_9_neigh_op_bot_5_49815),
    .O(seg_13_9_local_g1_5_53818)
  );
  LocalMux t2294 (
    .I(seg_13_9_neigh_op_bot_7_49817),
    .O(seg_13_9_local_g1_7_53820)
  );
  LocalMux t2295 (
    .I(seg_14_8_sp4_h_r_25_49946),
    .O(seg_14_8_local_g2_1_57529)
  );
  LocalMux t2296 (
    .I(seg_13_8_neigh_op_top_0_49933),
    .O(seg_13_8_local_g1_0_53690)
  );
  LocalMux t2297 (
    .I(seg_14_8_neigh_op_tnl_0_49933),
    .O(seg_14_8_local_g3_0_57536)
  );
  LocalMux t2298 (
    .I(seg_14_9_neigh_op_lft_0_49933),
    .O(seg_14_9_local_g0_0_57635)
  );
  LocalMux t2299 (
    .I(seg_13_8_neigh_op_top_1_49934),
    .O(seg_13_8_local_g0_1_53683)
  );
  CascadeMux t23 (
    .I(net_17292),
    .O(net_17292_cascademuxed)
  );
  CascadeMux t230 (
    .I(net_46700),
    .O(net_46700_cascademuxed)
  );
  LocalMux t2300 (
    .I(seg_13_9_lutff_1_out_49934),
    .O(seg_13_9_local_g1_1_53814)
  );
  LocalMux t2301 (
    .I(seg_14_9_neigh_op_lft_1_49934),
    .O(seg_14_9_local_g0_1_57636)
  );
  LocalMux t2302 (
    .I(seg_13_8_neigh_op_top_5_49938),
    .O(seg_13_8_local_g0_5_53687)
  );
  LocalMux t2303 (
    .I(seg_14_8_neigh_op_tnl_5_49938),
    .O(seg_14_8_local_g3_5_57541)
  );
  LocalMux t2304 (
    .I(seg_14_9_neigh_op_lft_5_49938),
    .O(seg_14_9_local_g0_5_57640)
  );
  LocalMux t2305 (
    .I(seg_13_8_neigh_op_top_6_49939),
    .O(seg_13_8_local_g0_6_53688)
  );
  LocalMux t2306 (
    .I(seg_13_9_lutff_6_out_49939),
    .O(seg_13_9_local_g2_6_53827)
  );
  LocalMux t2307 (
    .I(seg_14_9_neigh_op_lft_6_49939),
    .O(seg_14_9_local_g0_6_57641)
  );
  LocalMux t2308 (
    .I(seg_18_10_sp4_h_r_4_73181),
    .O(seg_18_10_local_g0_4_73085)
  );
  Span4Mux_h4 t2309 (
    .I(seg_18_10_sp4_h_l_45_57862),
    .O(seg_18_10_sp4_h_r_4_73181)
  );
  CascadeMux t231 (
    .I(net_46706),
    .O(net_46706_cascademuxed)
  );
  Span4Mux_h4 t2310 (
    .I(seg_14_10_sp4_v_b_8_53674),
    .O(seg_18_10_sp4_h_l_45_57862)
  );
  LocalMux t2311 (
    .I(seg_20_10_sp4_h_r_35_73178),
    .O(seg_20_10_local_g3_3_80139)
  );
  Span4Mux_h4 t2312 (
    .I(seg_18_10_sp4_h_l_45_57862),
    .O(seg_20_10_sp4_h_r_35_73178)
  );
  LocalMux t2313 (
    .I(seg_12_12_neigh_op_bnr_1_50180),
    .O(seg_12_12_local_g0_1_50344)
  );
  LocalMux t2314 (
    .I(seg_13_11_lutff_6_out_50185),
    .O(seg_13_11_local_g3_6_54081)
  );
  LocalMux t2315 (
    .I(seg_14_11_neigh_op_lft_6_50185),
    .O(seg_14_11_local_g0_6_57887)
  );
  LocalMux t2316 (
    .I(seg_14_13_neigh_op_bnl_1_50303),
    .O(seg_14_13_local_g3_1_58152)
  );
  LocalMux t2317 (
    .I(seg_13_13_neigh_op_bot_2_50304),
    .O(seg_13_13_local_g0_2_54299)
  );
  LocalMux t2318 (
    .I(seg_12_12_neigh_op_rgt_4_50306),
    .O(seg_12_12_local_g3_4_50371)
  );
  LocalMux t2319 (
    .I(seg_13_12_lutff_5_out_50307),
    .O(seg_13_12_local_g0_5_54179)
  );
  CascadeMux t232 (
    .I(net_46712),
    .O(net_46712_cascademuxed)
  );
  LocalMux t2320 (
    .I(seg_16_15_sp4_r_v_b_13_65895),
    .O(seg_16_15_local_g2_5_66055)
  );
  Span4Mux_v4 t2321 (
    .I(seg_17_12_sp4_h_l_37_54268),
    .O(seg_16_15_sp4_r_v_b_13_65895)
  );
  LocalMux t2322 (
    .I(seg_16_12_sp4_h_r_18_61937),
    .O(seg_16_12_local_g0_2_65667)
  );
  Span4Mux_h4 t2323 (
    .I(seg_15_12_sp4_h_l_41_46612),
    .O(seg_16_12_sp4_h_r_18_61937)
  );
  LocalMux t2324 (
    .I(seg_10_12_sp4_h_r_11_42778),
    .O(seg_10_12_local_g0_3_42684)
  );
  LocalMux t2325 (
    .I(seg_16_12_sp4_h_r_43_54276),
    .O(seg_16_12_local_g2_3_65684)
  );
  LocalMux t2326 (
    .I(seg_14_13_neigh_op_lft_3_50428),
    .O(seg_14_13_local_g0_3_58130)
  );
  LocalMux t2327 (
    .I(seg_13_12_neigh_op_top_4_50429),
    .O(seg_13_12_local_g0_4_54178)
  );
  LocalMux t2328 (
    .I(seg_13_13_lutff_4_out_50429),
    .O(seg_13_13_local_g3_4_54325)
  );
  LocalMux t2329 (
    .I(seg_13_13_lutff_5_out_50430),
    .O(seg_13_13_local_g2_5_54318)
  );
  CascadeMux t233 (
    .I(net_46805),
    .O(net_46805_cascademuxed)
  );
  LocalMux t2330 (
    .I(seg_13_14_neigh_op_bot_5_50430),
    .O(seg_13_14_local_g1_5_54433)
  );
  LocalMux t2331 (
    .I(seg_13_14_neigh_op_bot_6_50431),
    .O(seg_13_14_local_g0_6_54426)
  );
  LocalMux t2332 (
    .I(seg_18_13_sp4_h_r_29_65889),
    .O(seg_18_13_local_g3_5_73479)
  );
  Span4Mux_h4 t2333 (
    .I(seg_16_13_sp4_h_l_40_50567),
    .O(seg_18_13_sp4_h_r_29_65889)
  );
  LocalMux t2334 (
    .I(seg_10_13_sp4_h_r_23_39069),
    .O(seg_10_13_local_g0_7_42811)
  );
  Span4Mux_h4 t2335 (
    .I(seg_13_13_sp4_h_r_2_54395),
    .O(seg_10_13_sp4_h_r_23_39069)
  );
  LocalMux t2336 (
    .I(seg_16_13_sp4_h_r_19_62059),
    .O(seg_16_13_local_g0_3_65791)
  );
  Span4Mux_h4 t2337 (
    .I(seg_15_13_sp4_h_l_43_46737),
    .O(seg_16_13_sp4_h_r_19_62059)
  );
  LocalMux t2338 (
    .I(seg_15_13_sp4_h_r_28_54397),
    .O(seg_15_13_local_g2_4_61977)
  );
  LocalMux t2339 (
    .I(seg_11_13_sp4_h_r_20_42909),
    .O(seg_11_13_local_g1_4_46647)
  );
  CascadeMux t234 (
    .I(net_46823),
    .O(net_46823_cascademuxed)
  );
  LocalMux t2340 (
    .I(seg_19_14_sp4_h_r_17_73673),
    .O(seg_19_14_local_g0_1_77130)
  );
  Span4Mux_h4 t2341 (
    .I(seg_18_14_sp4_h_l_41_58350),
    .O(seg_19_14_sp4_h_r_17_73673)
  );
  Span4Mux_h4 t2342 (
    .I(seg_14_14_sp4_v_b_4_54162),
    .O(seg_18_14_sp4_h_l_41_58350)
  );
  LocalMux t2343 (
    .I(seg_12_13_neigh_op_tnr_2_50550),
    .O(seg_12_13_local_g3_2_50492)
  );
  LocalMux t2344 (
    .I(seg_14_14_neigh_op_lft_3_50551),
    .O(seg_14_14_local_g1_3_58261)
  );
  LocalMux t2345 (
    .I(seg_13_13_neigh_op_top_4_50552),
    .O(seg_13_13_local_g1_4_54309)
  );
  LocalMux t2346 (
    .I(seg_13_14_lutff_5_out_50553),
    .O(seg_13_14_local_g3_5_54449)
  );
  LocalMux t2347 (
    .I(seg_12_14_neigh_op_rgt_7_50555),
    .O(seg_12_14_local_g3_7_50620)
  );
  LocalMux t2348 (
    .I(seg_13_14_lutff_7_out_50555),
    .O(seg_13_14_local_g3_7_54451)
  );
  LocalMux t2349 (
    .I(seg_17_14_sp4_h_r_3_69841),
    .O(seg_17_14_local_g1_3_69753)
  );
  CascadeMux t235 (
    .I(net_46829),
    .O(net_46829_cascademuxed)
  );
  Span4Mux_h4 t2350 (
    .I(seg_17_14_sp4_h_l_37_54514),
    .O(seg_17_14_sp4_h_r_3_69841)
  );
  LocalMux t2351 (
    .I(seg_15_15_sp4_h_r_13_58467),
    .O(seg_15_15_local_g0_5_62208)
  );
  Span4Mux_h4 t2352 (
    .I(seg_14_15_sp4_v_b_0_54281),
    .O(seg_15_15_sp4_h_r_13_58467)
  );
  LocalMux t2353 (
    .I(seg_14_12_sp4_v_b_27_54159),
    .O(seg_14_12_local_g2_3_58023)
  );
  LocalMux t2354 (
    .I(seg_13_15_lutff_1_out_50672),
    .O(seg_13_15_local_g2_1_54560)
  );
  LocalMux t2355 (
    .I(seg_13_15_lutff_2_out_50673),
    .O(seg_13_15_local_g0_2_54545)
  );
  LocalMux t2356 (
    .I(seg_13_15_lutff_2_out_50673),
    .O(seg_13_15_local_g1_2_54553)
  );
  LocalMux t2357 (
    .I(seg_13_16_neigh_op_bot_4_50675),
    .O(seg_13_16_local_g0_4_54670)
  );
  LocalMux t2358 (
    .I(seg_13_16_neigh_op_bot_6_50677),
    .O(seg_13_16_local_g1_6_54680)
  );
  LocalMux t2359 (
    .I(seg_18_15_sp4_h_r_13_69959),
    .O(seg_18_15_local_g0_5_73701)
  );
  CascadeMux t236 (
    .I(net_46835),
    .O(net_46835_cascademuxed)
  );
  Span4Mux_h4 t2360 (
    .I(seg_17_15_sp4_h_l_37_54637),
    .O(seg_18_15_sp4_h_r_13_69959)
  );
  LocalMux t2361 (
    .I(seg_18_15_sp4_h_r_27_66133),
    .O(seg_18_15_local_g3_3_73723)
  );
  Span4Mux_h4 t2362 (
    .I(seg_16_15_sp4_h_l_38_50811),
    .O(seg_18_15_sp4_h_r_27_66133)
  );
  LocalMux t2363 (
    .I(seg_19_15_sp4_h_r_38_66133),
    .O(seg_19_15_local_g3_6_77261)
  );
  Span4Mux_h4 t2364 (
    .I(seg_16_15_sp4_h_l_38_50811),
    .O(seg_19_15_sp4_h_r_38_66133)
  );
  LocalMux t2365 (
    .I(seg_19_15_sp4_h_r_45_66138),
    .O(seg_19_15_local_g3_5_77260)
  );
  Span4Mux_h4 t2366 (
    .I(seg_16_15_sp4_h_l_40_50813),
    .O(seg_19_15_sp4_h_r_45_66138)
  );
  LocalMux t2367 (
    .I(seg_15_15_sp4_h_r_26_54641),
    .O(seg_15_15_local_g3_2_62229)
  );
  LocalMux t2368 (
    .I(seg_15_12_sp4_v_b_45_58119),
    .O(seg_15_12_local_g2_5_61855)
  );
  Span4Mux_v4 t2369 (
    .I(seg_15_15_sp4_h_l_39_46979),
    .O(seg_15_12_sp4_v_b_45_58119)
  );
  CascadeMux t237 (
    .I(net_46940),
    .O(net_46940_cascademuxed)
  );
  LocalMux t2370 (
    .I(seg_14_13_sp4_v_b_47_54414),
    .O(seg_14_13_local_g3_7_58158)
  );
  LocalMux t2371 (
    .I(seg_14_15_neigh_op_tnl_1_50795),
    .O(seg_14_15_local_g3_1_58398)
  );
  LocalMux t2372 (
    .I(seg_15_13_sp4_v_b_45_58242),
    .O(seg_15_13_local_g3_5_61986)
  );
  Span4Mux_v4 t2373 (
    .I(seg_15_16_sp4_h_l_39_47102),
    .O(seg_15_13_sp4_v_b_45_58242)
  );
  LocalMux t2374 (
    .I(seg_16_13_sp4_h_r_24_58221),
    .O(seg_16_13_local_g3_0_65812)
  );
  Span4Mux_h4 t2375 (
    .I(seg_14_13_sp4_v_t_37_54527),
    .O(seg_16_13_sp4_h_r_24_58221)
  );
  LocalMux t2376 (
    .I(seg_16_15_sp4_h_r_28_58473),
    .O(seg_16_15_local_g2_4_66054)
  );
  Span4Mux_h4 t2377 (
    .I(seg_14_15_sp4_v_t_41_54777),
    .O(seg_16_15_sp4_h_r_28_58473)
  );
  LocalMux t2378 (
    .I(seg_14_13_sp4_v_b_40_54407),
    .O(seg_14_13_local_g3_0_58151)
  );
  LocalMux t2379 (
    .I(seg_13_14_sp4_r_v_b_31_54409),
    .O(seg_13_14_local_g0_7_54427)
  );
  CascadeMux t238 (
    .I(net_47069),
    .O(net_47069_cascademuxed)
  );
  LocalMux t2380 (
    .I(seg_13_14_sp4_v_b_38_50697),
    .O(seg_13_14_local_g3_6_54450)
  );
  LocalMux t2381 (
    .I(seg_14_16_neigh_op_tnl_6_50923),
    .O(seg_14_16_local_g2_6_58518)
  );
  LocalMux t2382 (
    .I(seg_15_16_sp4_r_v_b_22_62196),
    .O(seg_15_16_local_g3_6_62356)
  );
  Span4Mux_v4 t2383 (
    .I(seg_16_17_sp4_h_l_40_51059),
    .O(seg_15_16_sp4_r_v_b_22_62196)
  );
  LocalMux t2384 (
    .I(seg_15_16_sp4_r_v_b_20_62194),
    .O(seg_15_16_local_g3_4_62354)
  );
  Span4Mux_v4 t2385 (
    .I(seg_16_17_sp4_h_l_44_51063),
    .O(seg_15_16_sp4_r_v_b_20_62194)
  );
  LocalMux t2386 (
    .I(seg_16_14_sp4_v_b_40_62190),
    .O(seg_16_14_local_g3_0_65935)
  );
  Span4Mux_v4 t2387 (
    .I(seg_16_17_sp4_h_l_46_51055),
    .O(seg_16_14_sp4_v_b_40_62190)
  );
  LocalMux t2388 (
    .I(seg_14_14_sp4_v_b_46_54536),
    .O(seg_14_14_local_g3_6_58280)
  );
  LocalMux t2389 (
    .I(seg_14_15_sp4_v_b_39_54652),
    .O(seg_14_15_local_g3_7_58404)
  );
  CascadeMux t239 (
    .I(net_47168),
    .O(net_47168_cascademuxed)
  );
  LocalMux t2390 (
    .I(seg_15_16_sp4_h_r_17_58596),
    .O(seg_15_16_local_g0_1_62327)
  );
  Span4Mux_h4 t2391 (
    .I(seg_14_16_sp4_v_t_41_54900),
    .O(seg_15_16_sp4_h_r_17_58596)
  );
  LocalMux t2392 (
    .I(seg_13_15_sp4_v_b_26_50698),
    .O(seg_13_15_local_g3_2_54569)
  );
  LocalMux t2393 (
    .I(seg_14_18_neigh_op_lft_3_51043),
    .O(seg_14_18_local_g0_3_58745)
  );
  LocalMux t2394 (
    .I(seg_12_18_neigh_op_rgt_4_51044),
    .O(seg_12_18_local_g2_4_51101)
  );
  LocalMux t2395 (
    .I(seg_14_18_neigh_op_lft_5_51045),
    .O(seg_14_18_local_g0_5_58747)
  );
  LocalMux t2396 (
    .I(seg_13_19_lutff_2_out_51165),
    .O(seg_13_19_local_g2_2_55053)
  );
  LocalMux t2397 (
    .I(seg_13_19_lutff_6_out_51169),
    .O(seg_13_19_local_g1_6_55049)
  );
  LocalMux t2398 (
    .I(seg_13_19_lutff_7_out_51170),
    .O(seg_13_19_local_g1_7_55050)
  );
  LocalMux t2399 (
    .I(seg_19_18_sp4_r_v_b_20_77427),
    .O(seg_19_18_local_g3_4_77565)
  );
  CascadeMux t24 (
    .I(net_17298),
    .O(net_17298_cascademuxed)
  );
  CascadeMux t240 (
    .I(net_47291),
    .O(net_47291_cascademuxed)
  );
  Span4Mux_v4 t2400 (
    .I(seg_20_19_sp4_h_l_38_66625),
    .O(seg_19_18_sp4_r_v_b_20_77427)
  );
  Span4Mux_h4 t2401 (
    .I(seg_16_19_sp4_h_l_42_51307),
    .O(seg_20_19_sp4_h_l_38_66625)
  );
  LocalMux t2402 (
    .I(seg_17_18_sp4_v_b_21_66272),
    .O(seg_17_18_local_g0_5_70239)
  );
  Span4Mux_v4 t2403 (
    .I(seg_17_19_sp4_h_l_39_55133),
    .O(seg_17_18_sp4_v_b_21_66272)
  );
  LocalMux t2404 (
    .I(seg_20_19_sp4_h_r_41_70457),
    .O(seg_20_19_local_g2_1_81236)
  );
  Span4Mux_h4 t2405 (
    .I(seg_17_19_sp4_h_l_45_55139),
    .O(seg_20_19_sp4_h_r_41_70457)
  );
  LocalMux t2406 (
    .I(seg_19_17_sp4_h_r_12_74037),
    .O(seg_19_17_local_g0_4_77439)
  );
  Span4Mux_h4 t2407 (
    .I(seg_18_17_sp4_h_l_36_58714),
    .O(seg_19_17_sp4_h_r_12_74037)
  );
  Span4Mux_h4 t2408 (
    .I(seg_14_17_sp4_v_t_36_55018),
    .O(seg_18_17_sp4_h_l_36_58714)
  );
  LocalMux t2409 (
    .I(seg_13_19_neigh_op_top_0_51286),
    .O(seg_13_19_local_g1_0_55043)
  );
  CascadeMux t241 (
    .I(net_47297),
    .O(net_47297_cascademuxed)
  );
  LocalMux t2410 (
    .I(seg_13_20_lutff_1_out_51287),
    .O(seg_13_20_local_g2_1_55175)
  );
  LocalMux t2411 (
    .I(seg_14_20_neigh_op_lft_4_51290),
    .O(seg_14_20_local_g0_4_58992)
  );
  LocalMux t2412 (
    .I(seg_13_20_lutff_5_out_51291),
    .O(seg_13_20_local_g1_5_55171)
  );
  LocalMux t2413 (
    .I(seg_14_20_neigh_op_lft_6_51292),
    .O(seg_14_20_local_g0_6_58994)
  );
  LocalMux t2414 (
    .I(seg_13_19_neigh_op_top_7_51293),
    .O(seg_13_19_local_g0_7_55042)
  );
  LocalMux t2415 (
    .I(seg_12_14_sp4_r_v_b_30_50579),
    .O(seg_12_14_local_g1_6_50603)
  );
  Span4Mux_v4 t2416 (
    .I(seg_13_16_sp4_v_t_43_51071),
    .O(seg_12_14_sp4_r_v_b_30_50579)
  );
  LocalMux t2417 (
    .I(seg_13_14_sp4_v_b_30_50579),
    .O(seg_13_14_local_g2_6_54442)
  );
  Span4Mux_v4 t2418 (
    .I(seg_13_16_sp4_v_t_43_51071),
    .O(seg_13_14_sp4_v_b_30_50579)
  );
  LocalMux t2419 (
    .I(seg_13_22_neigh_op_bot_6_51415),
    .O(seg_13_22_local_g1_6_55418)
  );
  CascadeMux t242 (
    .I(net_47420),
    .O(net_47420_cascademuxed)
  );
  LocalMux t2420 (
    .I(seg_12_12_sp4_r_v_b_33_50334),
    .O(seg_12_12_local_g2_1_50360)
  );
  Span4Mux_v4 t2421 (
    .I(seg_13_14_sp4_v_t_44_50826),
    .O(seg_12_12_sp4_r_v_b_33_50334)
  );
  Span4Mux_v4 t2422 (
    .I(seg_13_18_sp4_v_t_36_51310),
    .O(seg_13_14_sp4_v_t_44_50826)
  );
  LocalMux t2423 (
    .I(seg_12_14_sp4_r_v_b_5_50330),
    .O(seg_12_14_local_g1_5_50602)
  );
  Span4Mux_v4 t2424 (
    .I(seg_13_14_sp4_v_t_44_50826),
    .O(seg_12_14_sp4_r_v_b_5_50330)
  );
  LocalMux t2425 (
    .I(seg_13_22_lutff_1_out_51533),
    .O(seg_13_22_local_g0_1_55405)
  );
  LocalMux t2426 (
    .I(seg_12_21_neigh_op_tnr_3_51535),
    .O(seg_12_21_local_g3_3_51477)
  );
  LocalMux t2427 (
    .I(seg_13_22_lutff_5_out_51537),
    .O(seg_13_22_local_g1_5_55417)
  );
  LocalMux t2428 (
    .I(seg_12_21_neigh_op_tnr_7_51539),
    .O(seg_12_21_local_g2_7_51473)
  );
  LocalMux t2429 (
    .I(seg_12_21_sp4_h_r_44_40062),
    .O(seg_12_21_local_g2_4_51470)
  );
  CascadeMux t243 (
    .I(net_47543),
    .O(net_47543_cascademuxed)
  );
  Span4Mux_h4 t2430 (
    .I(seg_13_21_sp4_v_t_38_51681),
    .O(seg_12_21_sp4_h_r_44_40062)
  );
  LocalMux t2431 (
    .I(seg_13_27_lutff_2_out_52149),
    .O(seg_13_27_local_g2_2_56037)
  );
  LocalMux t2432 (
    .I(seg_12_27_neigh_op_rgt_4_52151),
    .O(seg_12_27_local_g2_4_52208)
  );
  LocalMux t2433 (
    .I(seg_13_27_lutff_4_out_52151),
    .O(seg_13_27_local_g3_4_56047)
  );
  LocalMux t2434 (
    .I(seg_12_27_neigh_op_rgt_5_52152),
    .O(seg_12_27_local_g2_5_52209)
  );
  LocalMux t2435 (
    .I(seg_13_27_lutff_5_out_52152),
    .O(seg_13_27_local_g2_5_56040)
  );
  LocalMux t2436 (
    .I(seg_14_27_neigh_op_lft_5_52152),
    .O(seg_14_27_local_g1_5_59862)
  );
  LocalMux t2437 (
    .I(seg_12_27_neigh_op_rgt_7_52154),
    .O(seg_12_27_local_g2_7_52211)
  );
  LocalMux t2438 (
    .I(seg_13_27_lutff_7_out_52154),
    .O(seg_13_27_local_g0_7_56026)
  );
  LocalMux t2439 (
    .I(seg_16_28_sp4_h_r_24_60066),
    .O(seg_16_28_local_g2_0_67649)
  );
  CascadeMux t244 (
    .I(net_47936),
    .O(net_47936_cascademuxed)
  );
  Span4Mux_h4 t2440 (
    .I(seg_14_28_sp4_v_b_0_55880),
    .O(seg_16_28_sp4_h_r_24_60066)
  );
  LocalMux t2441 (
    .I(seg_13_20_sp12_v_b_23_55128),
    .O(seg_13_20_local_g3_7_55189)
  );
  LocalMux t2442 (
    .I(seg_13_21_sp12_v_b_20_55128),
    .O(seg_13_21_local_g3_4_55309)
  );
  LocalMux t2443 (
    .I(seg_13_22_sp12_v_b_19_55128),
    .O(seg_13_22_local_g2_3_55423)
  );
  LocalMux t2444 (
    .I(seg_13_22_sp12_v_b_21_55250),
    .O(seg_13_22_local_g3_5_55433)
  );
  LocalMux t2445 (
    .I(seg_14_2_lutff_2_out_52869),
    .O(seg_14_2_local_g0_2_56776)
  );
  LocalMux t2446 (
    .I(seg_14_2_lutff_3_out_52870),
    .O(seg_14_2_local_g0_3_56777)
  );
  LocalMux t2447 (
    .I(seg_14_3_sp12_v_b_11_56584),
    .O(seg_14_3_local_g3_3_56924)
  );
  LocalMux t2448 (
    .I(seg_18_0_span4_vert_17_68222),
    .O(seg_18_0_local_g1_1_71885)
  );
  Span4Mux_v4 t2449 (
    .I(seg_18_2_sp4_h_l_47_56870),
    .O(seg_18_0_span4_vert_17_68222)
  );
  LocalMux t2450 (
    .I(seg_13_4_neigh_op_bnr_0_53026),
    .O(seg_13_4_local_g1_0_53198)
  );
  LocalMux t2451 (
    .I(seg_14_3_lutff_0_out_53026),
    .O(seg_14_3_local_g3_0_56921)
  );
  LocalMux t2452 (
    .I(seg_14_4_neigh_op_bot_0_53026),
    .O(seg_14_4_local_g1_0_57028)
  );
  LocalMux t2453 (
    .I(seg_14_3_lutff_1_out_53027),
    .O(seg_14_3_local_g2_1_56914)
  );
  LocalMux t2454 (
    .I(seg_14_3_lutff_2_out_53028),
    .O(seg_14_3_local_g0_2_56899)
  );
  LocalMux t2455 (
    .I(seg_14_2_neigh_op_top_3_53029),
    .O(seg_14_2_local_g1_3_56785)
  );
  LocalMux t2456 (
    .I(seg_15_3_neigh_op_lft_4_53030),
    .O(seg_15_3_local_g1_4_60739)
  );
  LocalMux t2457 (
    .I(seg_15_3_neigh_op_lft_5_53031),
    .O(seg_15_3_local_g0_5_60732)
  );
  LocalMux t2458 (
    .I(seg_14_4_neigh_op_bot_6_53032),
    .O(seg_14_4_local_g1_6_57034)
  );
  LocalMux t2459 (
    .I(seg_14_3_lutff_7_out_53033),
    .O(seg_14_3_local_g2_7_56920)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t246 (
    .carryinitin(),
    .carryinitout(t245)
  );
  LocalMux t2460 (
    .I(seg_13_4_neigh_op_rgt_0_53149),
    .O(seg_13_4_local_g3_0_53214)
  );
  LocalMux t2461 (
    .I(seg_14_3_neigh_op_top_0_53149),
    .O(seg_14_3_local_g0_0_56897)
  );
  LocalMux t2462 (
    .I(seg_14_4_lutff_0_out_53149),
    .O(seg_14_4_local_g3_0_57044)
  );
  LocalMux t2463 (
    .I(seg_13_3_neigh_op_tnr_1_53150),
    .O(seg_13_3_local_g3_1_53092)
  );
  LocalMux t2464 (
    .I(seg_13_4_neigh_op_rgt_1_53150),
    .O(seg_13_4_local_g3_1_53215)
  );
  LocalMux t2465 (
    .I(seg_14_3_neigh_op_top_1_53150),
    .O(seg_14_3_local_g1_1_56906)
  );
  LocalMux t2466 (
    .I(seg_13_4_neigh_op_rgt_2_53151),
    .O(seg_13_4_local_g2_2_53208)
  );
  LocalMux t2467 (
    .I(seg_14_4_lutff_2_out_53151),
    .O(seg_14_4_local_g2_2_57038)
  );
  LocalMux t2468 (
    .I(seg_13_3_neigh_op_tnr_4_53153),
    .O(seg_13_3_local_g3_4_53095)
  );
  LocalMux t2469 (
    .I(seg_13_4_neigh_op_rgt_4_53153),
    .O(seg_13_4_local_g2_4_53210)
  );
  LocalMux t2470 (
    .I(seg_14_3_neigh_op_top_4_53153),
    .O(seg_14_3_local_g1_4_56909)
  );
  LocalMux t2471 (
    .I(seg_14_4_lutff_5_out_53154),
    .O(seg_14_4_local_g3_5_57049)
  );
  LocalMux t2472 (
    .I(seg_13_4_neigh_op_rgt_7_53156),
    .O(seg_13_4_local_g3_7_53221)
  );
  LocalMux t2473 (
    .I(seg_14_3_neigh_op_top_7_53156),
    .O(seg_14_3_local_g0_7_56904)
  );
  LocalMux t2474 (
    .I(seg_14_4_lutff_7_out_53156),
    .O(seg_14_4_local_g0_7_57027)
  );
  LocalMux t2475 (
    .I(seg_14_4_lutff_7_out_53156),
    .O(seg_14_4_local_g3_7_57051)
  );
  LocalMux t2476 (
    .I(seg_14_7_lutff_1_out_53519),
    .O(seg_14_7_local_g3_1_57414)
  );
  LocalMux t2477 (
    .I(seg_13_8_neigh_op_bnr_6_53524),
    .O(seg_13_8_local_g1_6_53696)
  );
  LocalMux t2478 (
    .I(seg_14_7_lutff_6_out_53524),
    .O(seg_14_7_local_g1_6_57403)
  );
  LocalMux t2479 (
    .I(seg_14_8_neigh_op_bot_6_53524),
    .O(seg_14_8_local_g1_6_57526)
  );
  CascadeMux t248 (
    .I(net_48668),
    .O(net_48668_cascademuxed)
  );
  LocalMux t2480 (
    .I(seg_14_7_lutff_7_out_53525),
    .O(seg_14_7_local_g2_7_57412)
  );
  LocalMux t2481 (
    .I(seg_14_9_sp4_v_b_4_53547),
    .O(seg_14_9_local_g1_4_57647)
  );
  LocalMux t2482 (
    .I(seg_13_8_neigh_op_rgt_6_53647),
    .O(seg_13_8_local_g3_6_53712)
  );
  LocalMux t2483 (
    .I(seg_13_9_neigh_op_bnr_6_53647),
    .O(seg_13_9_local_g1_6_53819)
  );
  LocalMux t2484 (
    .I(seg_14_9_neigh_op_bot_6_53647),
    .O(seg_14_9_local_g1_6_57649)
  );
  LocalMux t2485 (
    .I(seg_13_8_neigh_op_rgt_7_53648),
    .O(seg_13_8_local_g3_7_53713)
  );
  LocalMux t2486 (
    .I(seg_14_8_lutff_7_out_53648),
    .O(seg_14_8_local_g1_7_57527)
  );
  LocalMux t2487 (
    .I(seg_14_9_neigh_op_bot_7_53648),
    .O(seg_14_9_local_g0_7_57642)
  );
  LocalMux t2488 (
    .I(seg_18_10_sp4_v_b_32_69242),
    .O(seg_18_10_local_g3_0_73105)
  );
  Span4Mux_v4 t2489 (
    .I(seg_18_8_sp4_h_l_45_57616),
    .O(seg_18_10_sp4_v_b_32_69242)
  );
  CascadeMux t249 (
    .I(net_48767),
    .O(net_48767_cascademuxed)
  );
  LocalMux t2490 (
    .I(seg_15_8_sp4_v_b_11_57259),
    .O(seg_15_8_local_g1_3_61353)
  );
  LocalMux t2491 (
    .I(seg_20_10_sp4_h_r_18_76804),
    .O(seg_20_10_local_g1_2_80122)
  );
  Span4Mux_h4 t2492 (
    .I(seg_19_10_sp4_h_l_42_61691),
    .O(seg_20_10_sp4_h_r_18_76804)
  );
  Span4Mux_h4 t2493 (
    .I(seg_15_10_sp4_v_b_1_57495),
    .O(seg_19_10_sp4_h_l_42_61691)
  );
  LocalMux t2494 (
    .I(seg_13_9_neigh_op_rgt_2_53766),
    .O(seg_13_9_local_g2_2_53823)
  );
  LocalMux t2495 (
    .I(seg_14_8_neigh_op_top_3_53767),
    .O(seg_14_8_local_g1_3_57523)
  );
  LocalMux t2496 (
    .I(seg_13_9_neigh_op_rgt_4_53768),
    .O(seg_13_9_local_g2_4_53825)
  );
  LocalMux t2497 (
    .I(seg_13_9_neigh_op_rgt_5_53769),
    .O(seg_13_9_local_g3_5_53834)
  );
  LocalMux t2498 (
    .I(seg_14_8_neigh_op_top_6_53770),
    .O(seg_14_8_local_g0_6_57518)
  );
  LocalMux t2499 (
    .I(seg_13_9_neigh_op_rgt_7_53771),
    .O(seg_13_9_local_g3_7_53836)
  );
  CascadeMux t25 (
    .I(net_17304),
    .O(net_17304_cascademuxed)
  );
  CascadeMux t250 (
    .I(net_48779),
    .O(net_48779_cascademuxed)
  );
  LocalMux t2500 (
    .I(seg_11_10_sp4_h_r_11_46363),
    .O(seg_11_10_local_g0_3_46269)
  );
  LocalMux t2501 (
    .I(seg_15_11_neigh_op_lft_0_54010),
    .O(seg_15_11_local_g1_0_61719)
  );
  LocalMux t2502 (
    .I(seg_14_11_lutff_1_out_54011),
    .O(seg_14_11_local_g1_1_57890)
  );
  LocalMux t2503 (
    .I(seg_14_11_lutff_3_out_54013),
    .O(seg_14_11_local_g0_3_57884)
  );
  LocalMux t2504 (
    .I(seg_14_12_neigh_op_bot_3_54013),
    .O(seg_14_12_local_g1_3_58015)
  );
  LocalMux t2505 (
    .I(seg_15_11_neigh_op_lft_5_54015),
    .O(seg_15_11_local_g0_5_61716)
  );
  LocalMux t2506 (
    .I(seg_15_11_neigh_op_lft_6_54016),
    .O(seg_15_11_local_g0_6_61717)
  );
  LocalMux t2507 (
    .I(seg_14_11_lutff_7_out_54017),
    .O(seg_14_11_local_g0_7_57888)
  );
  LocalMux t2508 (
    .I(seg_18_12_sp4_v_b_44_69610),
    .O(seg_18_12_local_g3_4_73355)
  );
  Span4Mux_v4 t2509 (
    .I(seg_18_11_sp4_h_l_41_57981),
    .O(seg_18_12_sp4_v_b_44_69610)
  );
  LocalMux t2510 (
    .I(seg_19_16_sp4_v_b_24_73803),
    .O(seg_19_16_local_g2_0_77349)
  );
  Span4Mux_v4 t2511 (
    .I(seg_19_14_sp4_h_l_37_62174),
    .O(seg_19_16_sp4_v_b_24_73803)
  );
  Span4Mux_h4 t2512 (
    .I(seg_15_14_sp4_v_b_0_57988),
    .O(seg_19_14_sp4_h_l_37_62174)
  );
  LocalMux t2513 (
    .I(seg_14_14_sp4_v_b_5_54161),
    .O(seg_14_14_local_g1_5_58263)
  );
  LocalMux t2514 (
    .I(seg_14_12_lutff_1_out_54134),
    .O(seg_14_12_local_g2_1_58021)
  );
  LocalMux t2515 (
    .I(seg_14_13_neigh_op_bot_2_54135),
    .O(seg_14_13_local_g1_2_58137)
  );
  LocalMux t2516 (
    .I(seg_14_13_neigh_op_bot_3_54136),
    .O(seg_14_13_local_g1_3_58138)
  );
  LocalMux t2517 (
    .I(seg_14_12_lutff_6_out_54139),
    .O(seg_14_12_local_g3_6_58034)
  );
  LocalMux t2518 (
    .I(seg_16_12_sp4_h_r_26_58102),
    .O(seg_16_12_local_g2_2_65683)
  );
  LocalMux t2519 (
    .I(seg_12_12_sp4_h_r_16_46613),
    .O(seg_12_12_local_g1_0_50351)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t252 (
    .carryinitin(),
    .carryinitout(t251)
  );
  LocalMux t2520 (
    .I(seg_12_12_sp4_h_r_18_46615),
    .O(seg_12_12_local_g1_2_50353)
  );
  LocalMux t2521 (
    .I(seg_18_13_sp4_h_r_39_62055),
    .O(seg_18_13_local_g2_7_73473)
  );
  Span4Mux_h4 t2522 (
    .I(seg_15_13_sp4_v_b_2_57867),
    .O(seg_18_13_sp4_h_r_39_62055)
  );
  LocalMux t2523 (
    .I(seg_19_14_sp4_h_r_4_77209),
    .O(seg_19_14_local_g1_4_77141)
  );
  Span4Mux_h4 t2524 (
    .I(seg_19_14_sp4_h_l_36_62175),
    .O(seg_19_14_sp4_h_r_4_77209)
  );
  Span4Mux_h4 t2525 (
    .I(seg_15_14_sp4_v_b_7_57993),
    .O(seg_19_14_sp4_h_l_36_62175)
  );
  LocalMux t2526 (
    .I(seg_18_13_sp4_r_v_b_20_73318),
    .O(seg_18_13_local_g3_4_73478)
  );
  Span4Mux_v4 t2527 (
    .I(seg_19_14_sp4_h_l_44_62185),
    .O(seg_18_13_sp4_r_v_b_20_73318)
  );
  Span4Mux_h4 t2528 (
    .I(seg_15_14_sp4_v_b_9_57995),
    .O(seg_19_14_sp4_h_l_44_62185)
  );
  LocalMux t2529 (
    .I(seg_19_14_sp4_h_r_5_77210),
    .O(seg_19_14_local_g0_5_77134)
  );
  Span4Mux_h4 t2530 (
    .I(seg_19_14_sp4_h_l_44_62185),
    .O(seg_19_14_sp4_h_r_5_77210)
  );
  LocalMux t2531 (
    .I(seg_15_14_neigh_op_bnl_2_54258),
    .O(seg_15_14_local_g2_2_62098)
  );
  LocalMux t2532 (
    .I(seg_14_13_lutff_7_out_54263),
    .O(seg_14_13_local_g1_7_58142)
  );
  LocalMux t2533 (
    .I(seg_22_13_sp4_h_r_9_88248),
    .O(seg_22_13_local_g1_1_88152)
  );
  Span4Mux_h4 t2534 (
    .I(seg_22_13_sp4_h_l_36_73545),
    .O(seg_22_13_sp4_h_r_9_88248)
  );
  Span4Mux_h4 t2535 (
    .I(seg_18_13_sp4_h_l_47_58223),
    .O(seg_22_13_sp4_h_l_36_73545)
  );
  LocalMux t2536 (
    .I(seg_16_13_sp4_h_r_26_58225),
    .O(seg_16_13_local_g2_2_65806)
  );
  LocalMux t2537 (
    .I(seg_19_13_sp4_h_r_16_73551),
    .O(seg_19_13_local_g1_0_77035)
  );
  Span4Mux_h4 t2538 (
    .I(seg_18_13_sp4_h_l_39_58225),
    .O(seg_19_13_sp4_h_r_16_73551)
  );
  LocalMux t2539 (
    .I(seg_19_13_sp4_h_r_38_65887),
    .O(seg_19_13_local_g2_6_77049)
  );
  Span4Mux_h4 t2540 (
    .I(seg_16_13_sp4_h_l_37_50560),
    .O(seg_19_13_sp4_h_r_38_65887)
  );
  LocalMux t2541 (
    .I(seg_19_13_sp4_h_r_47_65884),
    .O(seg_19_13_local_g2_7_77050)
  );
  Span4Mux_h4 t2542 (
    .I(seg_16_13_sp4_h_l_39_50564),
    .O(seg_19_13_sp4_h_r_47_65884)
  );
  LocalMux t2543 (
    .I(seg_14_13_sp4_h_r_30_50568),
    .O(seg_14_13_local_g3_6_58157)
  );
  LocalMux t2544 (
    .I(seg_12_13_sp4_h_r_8_50570),
    .O(seg_12_13_local_g1_0_50474)
  );
  LocalMux t2545 (
    .I(seg_18_12_sp4_v_b_19_69363),
    .O(seg_18_12_local_g0_3_73330)
  );
  Span4Mux_v4 t2546 (
    .I(seg_18_13_sp4_h_l_43_58229),
    .O(seg_18_12_sp4_v_b_19_69363)
  );
  LocalMux t2547 (
    .I(seg_18_13_sp4_h_r_11_73547),
    .O(seg_18_13_local_g1_3_73461)
  );
  Span4Mux_h4 t2548 (
    .I(seg_18_13_sp4_h_l_45_58231),
    .O(seg_18_13_sp4_h_r_11_73547)
  );
  LocalMux t2549 (
    .I(seg_19_16_sp4_h_r_5_77414),
    .O(seg_19_16_local_g1_5_77346)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t255 (
    .carryinitin(),
    .carryinitout(t254)
  );
  Span4Mux_h4 t2550 (
    .I(seg_19_16_sp4_h_l_39_62424),
    .O(seg_19_16_sp4_h_r_5_77414)
  );
  Span4Mux_h4 t2551 (
    .I(seg_15_16_sp4_v_b_2_58236),
    .O(seg_19_16_sp4_h_l_39_62424)
  );
  LocalMux t2552 (
    .I(seg_19_14_sp4_h_r_20_73678),
    .O(seg_19_14_local_g0_4_77133)
  );
  Span4Mux_h4 t2553 (
    .I(seg_18_14_sp4_h_l_36_58345),
    .O(seg_19_14_sp4_h_r_20_73678)
  );
  Span4Mux_h4 t2554 (
    .I(seg_14_14_sp4_v_b_1_54157),
    .O(seg_18_14_sp4_h_l_36_58345)
  );
  LocalMux t2555 (
    .I(seg_20_14_sp4_h_r_31_73676),
    .O(seg_20_14_local_g3_7_80635)
  );
  Span4Mux_h4 t2556 (
    .I(seg_18_14_sp4_h_l_42_58353),
    .O(seg_20_14_sp4_h_r_31_73676)
  );
  Span4Mux_h4 t2557 (
    .I(seg_14_14_sp4_v_b_1_54157),
    .O(seg_18_14_sp4_h_l_42_58353)
  );
  LocalMux t2558 (
    .I(seg_15_13_neigh_op_tnl_1_54380),
    .O(seg_15_13_local_g2_1_61974)
  );
  LocalMux t2559 (
    .I(seg_14_14_lutff_5_out_54384),
    .O(seg_14_14_local_g3_5_58279)
  );
  LocalMux t2560 (
    .I(seg_14_14_lutff_6_out_54385),
    .O(seg_14_14_local_g2_6_58272)
  );
  LocalMux t2561 (
    .I(seg_15_14_neigh_op_lft_6_54385),
    .O(seg_15_14_local_g0_6_62086)
  );
  LocalMux t2562 (
    .I(seg_18_15_sp4_v_b_37_69972),
    .O(seg_18_15_local_g3_5_73725)
  );
  Span4Mux_v4 t2563 (
    .I(seg_18_14_sp4_h_l_37_58344),
    .O(seg_18_15_sp4_v_b_37_69972)
  );
  LocalMux t2564 (
    .I(seg_17_14_sp4_h_r_6_69844),
    .O(seg_17_14_local_g1_6_69756)
  );
  Span4Mux_h4 t2565 (
    .I(seg_17_14_sp4_h_l_38_54519),
    .O(seg_17_14_sp4_h_r_6_69844)
  );
  LocalMux t2566 (
    .I(seg_17_14_sp4_h_r_0_69836),
    .O(seg_17_14_local_g1_0_69750)
  );
  Span4Mux_h4 t2567 (
    .I(seg_17_14_sp4_h_l_44_54525),
    .O(seg_17_14_sp4_h_r_0_69836)
  );
  LocalMux t2568 (
    .I(seg_15_12_sp4_v_b_47_58121),
    .O(seg_15_12_local_g2_7_61857)
  );
  LocalMux t2569 (
    .I(seg_19_16_sp4_h_r_9_77418),
    .O(seg_19_16_local_g0_1_77334)
  );
  CascadeMux t257 (
    .I(net_49892),
    .O(net_49892_cascademuxed)
  );
  Span4Mux_h4 t2570 (
    .I(seg_19_16_sp4_h_l_44_62431),
    .O(seg_19_16_sp4_h_r_9_77418)
  );
  Span4Mux_h4 t2571 (
    .I(seg_15_16_sp4_v_b_9_58241),
    .O(seg_19_16_sp4_h_l_44_62431)
  );
  LocalMux t2572 (
    .I(seg_19_15_sp4_h_r_16_73797),
    .O(seg_19_15_local_g1_0_77239)
  );
  Span4Mux_h4 t2573 (
    .I(seg_18_15_sp4_h_l_44_58478),
    .O(seg_19_15_sp4_h_r_16_73797)
  );
  Span4Mux_h4 t2574 (
    .I(seg_14_15_sp4_v_b_3_54282),
    .O(seg_18_15_sp4_h_l_44_58478)
  );
  LocalMux t2575 (
    .I(seg_19_15_sp4_h_r_19_73798),
    .O(seg_19_15_local_g0_3_77234)
  );
  Span4Mux_h4 t2576 (
    .I(seg_18_15_sp4_h_l_38_58472),
    .O(seg_19_15_sp4_h_r_19_73798)
  );
  Span4Mux_h4 t2577 (
    .I(seg_14_15_sp4_v_b_9_54288),
    .O(seg_18_15_sp4_h_l_38_58472)
  );
  LocalMux t2578 (
    .I(seg_14_11_sp4_v_b_45_54166),
    .O(seg_14_11_local_g2_5_57902)
  );
  LocalMux t2579 (
    .I(seg_14_14_neigh_op_top_0_54502),
    .O(seg_14_14_local_g1_0_58258)
  );
  CascadeMux t258 (
    .I(net_49922),
    .O(net_49922_cascademuxed)
  );
  LocalMux t2580 (
    .I(seg_14_16_neigh_op_bot_0_54502),
    .O(seg_14_16_local_g1_0_58504)
  );
  LocalMux t2581 (
    .I(seg_13_15_neigh_op_rgt_2_54504),
    .O(seg_13_15_local_g2_2_54561)
  );
  LocalMux t2582 (
    .I(seg_14_14_neigh_op_top_4_54506),
    .O(seg_14_14_local_g1_4_58262)
  );
  LocalMux t2583 (
    .I(seg_14_16_neigh_op_bot_4_54506),
    .O(seg_14_16_local_g0_4_58500)
  );
  LocalMux t2584 (
    .I(seg_13_15_neigh_op_rgt_6_54508),
    .O(seg_13_15_local_g3_6_54573)
  );
  LocalMux t2585 (
    .I(seg_14_15_lutff_6_out_54508),
    .O(seg_14_15_local_g1_6_58387)
  );
  LocalMux t2586 (
    .I(seg_14_16_neigh_op_bot_7_54509),
    .O(seg_14_16_local_g1_7_58511)
  );
  LocalMux t2587 (
    .I(seg_16_15_sp4_h_r_38_54642),
    .O(seg_16_15_local_g2_6_66056)
  );
  LocalMux t2588 (
    .I(seg_16_12_sp4_h_r_14_61933),
    .O(seg_16_12_local_g1_6_65679)
  );
  Span4Mux_h4 t2589 (
    .I(seg_15_12_sp4_v_t_47_58244),
    .O(seg_16_12_sp4_h_r_14_61933)
  );
  CascadeMux t259 (
    .I(net_50261),
    .O(net_50261_cascademuxed)
  );
  LocalMux t2590 (
    .I(seg_14_13_sp4_v_b_34_54291),
    .O(seg_14_13_local_g2_2_58145)
  );
  LocalMux t2591 (
    .I(seg_14_12_sp4_v_b_39_54283),
    .O(seg_14_12_local_g2_7_58027)
  );
  LocalMux t2592 (
    .I(seg_14_13_sp4_v_b_28_54285),
    .O(seg_14_13_local_g3_4_58155)
  );
  LocalMux t2593 (
    .I(seg_13_16_neigh_op_rgt_0_54625),
    .O(seg_13_16_local_g2_0_54682)
  );
  LocalMux t2594 (
    .I(seg_13_16_neigh_op_rgt_3_54628),
    .O(seg_13_16_local_g3_3_54693)
  );
  LocalMux t2595 (
    .I(seg_14_16_lutff_5_out_54630),
    .O(seg_14_16_local_g0_5_58501)
  );
  LocalMux t2596 (
    .I(seg_15_15_neigh_op_tnl_5_54630),
    .O(seg_15_15_local_g2_5_62224)
  );
  LocalMux t2597 (
    .I(seg_13_16_neigh_op_rgt_6_54631),
    .O(seg_13_16_local_g3_6_54696)
  );
  LocalMux t2598 (
    .I(seg_13_16_neigh_op_rgt_7_54632),
    .O(seg_13_16_local_g2_7_54689)
  );
  LocalMux t2599 (
    .I(seg_14_14_sp4_v_b_26_54406),
    .O(seg_14_14_local_g3_2_58276)
  );
  CascadeMux t26 (
    .I(net_17397),
    .O(net_17397_cascademuxed)
  );
  CascadeMux t260 (
    .I(net_50273),
    .O(net_50273_cascademuxed)
  );
  LocalMux t2600 (
    .I(seg_14_13_sp4_v_b_45_54412),
    .O(seg_14_13_local_g2_5_58148)
  );
  LocalMux t2601 (
    .I(seg_14_17_lutff_1_out_54749),
    .O(seg_14_17_local_g3_1_58644)
  );
  LocalMux t2602 (
    .I(seg_13_17_neigh_op_rgt_2_54750),
    .O(seg_13_17_local_g3_2_54815)
  );
  LocalMux t2603 (
    .I(seg_13_17_neigh_op_rgt_3_54751),
    .O(seg_13_17_local_g2_3_54808)
  );
  LocalMux t2604 (
    .I(seg_13_17_neigh_op_rgt_7_54755),
    .O(seg_13_17_local_g2_7_54812)
  );
  LocalMux t2605 (
    .I(seg_14_14_sp4_v_b_47_54537),
    .O(seg_14_14_local_g3_7_58281)
  );
  LocalMux t2606 (
    .I(seg_14_18_lutff_0_out_54871),
    .O(seg_14_18_local_g3_0_58766)
  );
  LocalMux t2607 (
    .I(seg_14_18_lutff_1_out_54872),
    .O(seg_14_18_local_g3_1_58767)
  );
  LocalMux t2608 (
    .I(seg_14_18_lutff_3_out_54874),
    .O(seg_14_18_local_g1_3_58753)
  );
  LocalMux t2609 (
    .I(seg_14_18_lutff_5_out_54876),
    .O(seg_14_18_local_g2_5_58763)
  );
  CascadeMux t261 (
    .I(net_50378),
    .O(net_50378_cascademuxed)
  );
  LocalMux t2610 (
    .I(seg_17_18_sp4_h_r_3_70333),
    .O(seg_17_18_local_g1_3_70245)
  );
  Span4Mux_h4 t2611 (
    .I(seg_17_18_sp4_h_l_38_55011),
    .O(seg_17_18_sp4_h_r_3_70333)
  );
  LocalMux t2612 (
    .I(seg_19_18_sp4_h_r_27_70333),
    .O(seg_19_18_local_g3_3_77564)
  );
  Span4Mux_h4 t2613 (
    .I(seg_17_18_sp4_h_l_38_55011),
    .O(seg_19_18_sp4_h_r_27_70333)
  );
  LocalMux t2614 (
    .I(seg_18_17_sp4_v_b_21_69980),
    .O(seg_18_17_local_g1_5_73955)
  );
  Span4Mux_v4 t2615 (
    .I(seg_18_18_sp4_h_l_45_58846),
    .O(seg_18_17_sp4_v_b_21_69980)
  );
  LocalMux t2616 (
    .I(seg_19_17_sp4_h_r_4_77515),
    .O(seg_19_17_local_g1_4_77447)
  );
  Span4Mux_h4 t2617 (
    .I(seg_19_17_sp4_h_l_41_62549),
    .O(seg_19_17_sp4_h_r_4_77515)
  );
  Span4Mux_h4 t2618 (
    .I(seg_15_17_sp4_v_t_41_58853),
    .O(seg_19_17_sp4_h_l_41_62549)
  );
  LocalMux t2619 (
    .I(seg_14_19_lutff_0_out_54994),
    .O(seg_14_19_local_g1_0_58873)
  );
  CascadeMux t262 (
    .I(net_50384),
    .O(net_50384_cascademuxed)
  );
  LocalMux t2620 (
    .I(seg_15_18_neigh_op_tnl_1_54995),
    .O(seg_15_18_local_g3_1_62597)
  );
  LocalMux t2621 (
    .I(seg_13_19_neigh_op_rgt_6_55000),
    .O(seg_13_19_local_g2_6_55057)
  );
  LocalMux t2622 (
    .I(seg_13_19_neigh_op_rgt_7_55001),
    .O(seg_13_19_local_g2_7_55058)
  );
  LocalMux t2623 (
    .I(seg_14_19_neigh_op_top_0_55117),
    .O(seg_14_19_local_g0_0_58865)
  );
  LocalMux t2624 (
    .I(seg_14_20_lutff_1_out_55118),
    .O(seg_14_20_local_g2_1_59005)
  );
  LocalMux t2625 (
    .I(seg_14_20_lutff_2_out_55119),
    .O(seg_14_20_local_g3_2_59014)
  );
  LocalMux t2626 (
    .I(seg_14_19_neigh_op_top_4_55121),
    .O(seg_14_19_local_g1_4_58877)
  );
  LocalMux t2627 (
    .I(seg_18_17_sp4_v_b_47_70228),
    .O(seg_18_17_local_g2_7_73965)
  );
  Span4Mux_v4 t2628 (
    .I(seg_18_20_sp4_h_l_47_59084),
    .O(seg_18_17_sp4_v_b_47_70228)
  );
  LocalMux t2629 (
    .I(seg_19_17_sp4_v_b_14_73804),
    .O(seg_19_17_local_g1_6_77449)
  );
  CascadeMux t263 (
    .I(net_50390),
    .O(net_50390_cascademuxed)
  );
  Span4Mux_v4 t2630 (
    .I(seg_19_18_sp4_h_l_38_62671),
    .O(seg_19_17_sp4_v_b_14_73804)
  );
  Span4Mux_h4 t2631 (
    .I(seg_15_18_sp4_v_t_38_58973),
    .O(seg_19_18_sp4_h_l_38_62671)
  );
  LocalMux t2632 (
    .I(seg_14_18_sp4_v_b_38_55020),
    .O(seg_14_18_local_g2_6_58764)
  );
  LocalMux t2633 (
    .I(seg_14_20_neigh_op_top_7_55247),
    .O(seg_14_20_local_g0_7_58995)
  );
  LocalMux t2634 (
    .I(seg_14_26_lutff_3_out_55858),
    .O(seg_14_26_local_g3_3_59753)
  );
  LocalMux t2635 (
    .I(seg_16_28_sp4_h_r_12_63897),
    .O(seg_16_28_local_g1_4_67645)
  );
  Span4Mux_h4 t2636 (
    .I(seg_15_28_sp4_v_b_1_59709),
    .O(seg_16_28_sp4_h_r_12_63897)
  );
  LocalMux t2637 (
    .I(seg_14_27_lutff_2_out_55980),
    .O(seg_14_27_local_g1_2_59859)
  );
  LocalMux t2638 (
    .I(seg_14_27_lutff_5_out_55983),
    .O(seg_14_27_local_g2_5_59870)
  );
  LocalMux t2639 (
    .I(seg_15_29_sp4_v_b_11_59842),
    .O(seg_15_29_local_g1_3_63936)
  );
  CascadeMux t264 (
    .I(net_50396),
    .O(net_50396_cascademuxed)
  );
  LocalMux t2640 (
    .I(seg_13_27_sp4_v_b_18_52054),
    .O(seg_13_27_local_g0_2_56021)
  );
  Span4Mux_v4 t2641 (
    .I(seg_13_28_sp4_h_r_7_56245),
    .O(seg_13_27_sp4_v_b_18_52054)
  );
  LocalMux t2642 (
    .I(seg_12_27_sp4_v_b_19_48224),
    .O(seg_12_27_local_g1_3_52199)
  );
  Span4Mux_v4 t2643 (
    .I(seg_12_28_sp4_h_l_43_37089),
    .O(seg_12_27_sp4_v_b_19_48224)
  );
  Span4Mux_h4 t2644 (
    .I(seg_12_28_sp4_h_r_10_52407),
    .O(seg_12_28_sp4_h_l_43_37089)
  );
  LocalMux t2645 (
    .I(seg_12_28_sp4_h_r_10_52407),
    .O(seg_12_28_local_g0_2_52313)
  );
  LocalMux t2646 (
    .I(seg_14_2_neigh_op_rgt_0_56697),
    .O(seg_14_2_local_g2_0_56790)
  );
  LocalMux t2647 (
    .I(seg_14_3_neigh_op_bnr_0_56697),
    .O(seg_14_3_local_g1_0_56905)
  );
  LocalMux t2648 (
    .I(seg_15_2_lutff_0_out_56697),
    .O(seg_15_2_local_g0_0_60604)
  );
  LocalMux t2649 (
    .I(seg_15_3_neigh_op_bot_0_56697),
    .O(seg_15_3_local_g1_0_60735)
  );
  CascadeMux t265 (
    .I(net_50402),
    .O(net_50402_cascademuxed)
  );
  LocalMux t2650 (
    .I(seg_16_2_neigh_op_lft_0_56697),
    .O(seg_16_2_local_g1_0_64443)
  );
  LocalMux t2651 (
    .I(seg_14_3_neigh_op_bnr_1_56698),
    .O(seg_14_3_local_g0_1_56898)
  );
  LocalMux t2652 (
    .I(seg_16_2_neigh_op_lft_1_56698),
    .O(seg_16_2_local_g0_1_64436)
  );
  LocalMux t2653 (
    .I(seg_15_2_lutff_2_out_56699),
    .O(seg_15_2_local_g0_2_60606)
  );
  LocalMux t2654 (
    .I(seg_15_3_neigh_op_bot_2_56699),
    .O(seg_15_3_local_g0_2_60729)
  );
  LocalMux t2655 (
    .I(seg_15_2_lutff_6_out_56703),
    .O(seg_15_2_local_g0_6_60610)
  );
  LocalMux t2656 (
    .I(seg_16_2_neigh_op_lft_6_56703),
    .O(seg_16_2_local_g1_6_64449)
  );
  LocalMux t2657 (
    .I(seg_17_0_span4_horz_r_11_60434),
    .O(seg_17_0_local_g1_3_68056)
  );
  IoSpan4Mux t2658 (
    .I(seg_15_0_span4_vert_19_56732),
    .O(seg_17_0_span4_horz_r_11_60434)
  );
  LocalMux t2659 (
    .I(seg_15_3_lutff_1_out_56857),
    .O(seg_15_3_local_g1_1_60736)
  );
  CascadeMux t266 (
    .I(net_50408),
    .O(net_50408_cascademuxed)
  );
  LocalMux t2660 (
    .I(seg_14_2_neigh_op_tnr_2_56858),
    .O(seg_14_2_local_g3_2_56800)
  );
  LocalMux t2661 (
    .I(seg_14_3_neigh_op_rgt_2_56858),
    .O(seg_14_3_local_g2_2_56915)
  );
  LocalMux t2662 (
    .I(seg_15_2_neigh_op_top_2_56858),
    .O(seg_15_2_local_g1_2_60614)
  );
  LocalMux t2663 (
    .I(seg_15_3_lutff_2_out_56858),
    .O(seg_15_3_local_g3_2_60753)
  );
  LocalMux t2664 (
    .I(seg_14_2_neigh_op_tnr_3_56859),
    .O(seg_14_2_local_g2_3_56793)
  );
  LocalMux t2665 (
    .I(seg_14_3_neigh_op_rgt_3_56859),
    .O(seg_14_3_local_g2_3_56916)
  );
  LocalMux t2666 (
    .I(seg_15_2_neigh_op_top_3_56859),
    .O(seg_15_2_local_g1_3_60615)
  );
  LocalMux t2667 (
    .I(seg_15_3_lutff_3_out_56859),
    .O(seg_15_3_local_g1_3_60738)
  );
  LocalMux t2668 (
    .I(seg_15_3_lutff_4_out_56860),
    .O(seg_15_3_local_g2_4_60747)
  );
  LocalMux t2669 (
    .I(seg_15_3_lutff_6_out_56862),
    .O(seg_15_3_local_g2_6_60749)
  );
  CascadeMux t267 (
    .I(net_50414),
    .O(net_50414_cascademuxed)
  );
  LocalMux t2670 (
    .I(seg_14_2_neigh_op_tnr_7_56863),
    .O(seg_14_2_local_g3_7_56805)
  );
  LocalMux t2671 (
    .I(seg_14_3_neigh_op_rgt_7_56863),
    .O(seg_14_3_local_g3_7_56928)
  );
  LocalMux t2672 (
    .I(seg_15_2_neigh_op_top_7_56863),
    .O(seg_15_2_local_g0_7_60611)
  );
  LocalMux t2673 (
    .I(seg_15_3_lutff_7_out_56863),
    .O(seg_15_3_local_g3_7_60758)
  );
  LocalMux t2674 (
    .I(seg_16_2_neigh_op_tnl_7_56863),
    .O(seg_16_2_local_g2_7_64458)
  );
  LocalMux t2675 (
    .I(seg_16_2_neigh_op_tnl_7_56863),
    .O(seg_16_2_local_g3_7_64466)
  );
  LocalMux t2676 (
    .I(seg_15_6_sp4_h_r_43_49707),
    .O(seg_15_6_local_g3_3_61123)
  );
  Span4Mux_h4 t2677 (
    .I(seg_16_6_sp4_v_b_6_60840),
    .O(seg_15_6_sp4_h_r_43_49707)
  );
  LocalMux t2678 (
    .I(seg_16_9_sp4_v_b_19_61332),
    .O(seg_16_9_local_g1_3_65307)
  );
  Span4Mux_v4 t2679 (
    .I(seg_16_6_sp4_h_l_36_49700),
    .O(seg_16_9_sp4_v_b_19_61332)
  );
  CascadeMux t268 (
    .I(net_50420),
    .O(net_50420_cascademuxed)
  );
  LocalMux t2680 (
    .I(seg_15_10_sp4_r_v_b_17_61453),
    .O(seg_15_10_local_g3_1_61613)
  );
  Span4Mux_v4 t2681 (
    .I(seg_16_7_sp4_v_b_8_60965),
    .O(seg_15_10_sp4_r_v_b_17_61453)
  );
  LocalMux t2682 (
    .I(seg_15_9_sp4_r_v_b_0_61203),
    .O(seg_15_9_local_g1_0_61473)
  );
  LocalMux t2683 (
    .I(seg_16_9_sp4_v_b_0_61203),
    .O(seg_16_9_local_g1_0_65304)
  );
  LocalMux t2684 (
    .I(seg_14_9_neigh_op_bnr_0_57471),
    .O(seg_14_9_local_g1_0_57643)
  );
  LocalMux t2685 (
    .I(seg_15_8_lutff_0_out_57471),
    .O(seg_15_8_local_g1_0_61350)
  );
  LocalMux t2686 (
    .I(seg_13_8_sp4_h_r_8_53786),
    .O(seg_13_8_local_g0_0_53682)
  );
  LocalMux t2687 (
    .I(seg_13_9_sp4_h_r_20_50079),
    .O(seg_13_9_local_g1_4_53817)
  );
  Span4Mux_h4 t2688 (
    .I(seg_16_9_sp4_v_b_4_61207),
    .O(seg_13_9_sp4_h_r_20_50079)
  );
  LocalMux t2689 (
    .I(seg_15_10_neigh_op_bot_0_57594),
    .O(seg_15_10_local_g1_0_61596)
  );
  CascadeMux t269 (
    .I(net_50501),
    .O(net_50501_cascademuxed)
  );
  LocalMux t2690 (
    .I(seg_14_10_neigh_op_bnr_5_57599),
    .O(seg_14_10_local_g0_5_57763)
  );
  LocalMux t2691 (
    .I(seg_15_10_neigh_op_bot_5_57599),
    .O(seg_15_10_local_g1_5_61601)
  );
  LocalMux t2692 (
    .I(seg_15_11_sp12_v_b_10_60942),
    .O(seg_15_11_local_g2_2_61729)
  );
  LocalMux t2693 (
    .I(seg_15_10_sp4_v_b_19_57625),
    .O(seg_15_10_local_g1_3_61599)
  );
  LocalMux t2694 (
    .I(seg_15_12_sp4_v_b_11_57751),
    .O(seg_15_12_local_g1_3_61845)
  );
  LocalMux t2695 (
    .I(seg_14_11_neigh_op_bnr_4_57721),
    .O(seg_14_11_local_g1_4_57893)
  );
  LocalMux t2696 (
    .I(seg_15_10_lutff_4_out_57721),
    .O(seg_15_10_local_g0_4_61592)
  );
  LocalMux t2697 (
    .I(seg_15_14_sp12_v_b_4_60943),
    .O(seg_15_14_local_g2_4_62100)
  );
  LocalMux t2698 (
    .I(seg_21_10_sp4_h_r_37_73175),
    .O(seg_21_10_local_g2_5_83964)
  );
  Span4Mux_h4 t2699 (
    .I(seg_18_10_sp4_h_l_44_57863),
    .O(seg_21_10_sp4_h_r_37_73175)
  );
  CascadeMux t27 (
    .I(net_17415),
    .O(net_17415_cascademuxed)
  );
  CascadeMux t270 (
    .I(net_50507),
    .O(net_50507_cascademuxed)
  );
  LocalMux t2700 (
    .I(seg_12_18_sp4_r_v_b_6_50825),
    .O(seg_12_18_local_g1_6_51095)
  );
  Span4Mux_v4 t2701 (
    .I(seg_13_14_sp4_v_b_6_50333),
    .O(seg_12_18_sp4_r_v_b_6_50825)
  );
  Span4Mux_v4 t2702 (
    .I(seg_13_10_sp4_h_r_0_54022),
    .O(seg_13_14_sp4_v_b_6_50333)
  );
  LocalMux t2703 (
    .I(seg_13_13_sp4_v_b_19_50333),
    .O(seg_13_13_local_g0_3_54300)
  );
  Span4Mux_v4 t2704 (
    .I(seg_13_10_sp4_h_r_0_54022),
    .O(seg_13_13_sp4_v_b_19_50333)
  );
  LocalMux t2705 (
    .I(seg_13_15_sp4_v_b_43_50825),
    .O(seg_13_15_local_g3_3_54570)
  );
  Span4Mux_v4 t2706 (
    .I(seg_13_14_sp4_v_b_6_50333),
    .O(seg_13_15_sp4_v_b_43_50825)
  );
  LocalMux t2707 (
    .I(seg_13_19_sp4_v_b_44_51318),
    .O(seg_13_19_local_g2_4_55055)
  );
  Span4Mux_v4 t2708 (
    .I(seg_13_18_sp4_v_b_6_50825),
    .O(seg_13_19_sp4_v_b_44_51318)
  );
  Span4Mux_v4 t2709 (
    .I(seg_13_14_sp4_v_b_6_50333),
    .O(seg_13_18_sp4_v_b_6_50825)
  );
  CascadeMux t271 (
    .I(net_50513),
    .O(net_50513_cascademuxed)
  );
  LocalMux t2710 (
    .I(seg_13_19_sp4_v_b_44_51318),
    .O(seg_13_19_local_g3_4_55063)
  );
  LocalMux t2711 (
    .I(seg_17_12_sp4_v_b_29_65652),
    .O(seg_17_12_local_g3_5_69525)
  );
  Span4Mux_v4 t2712 (
    .I(seg_17_10_sp4_h_l_37_54022),
    .O(seg_17_12_sp4_v_b_29_65652)
  );
  LocalMux t2713 (
    .I(seg_17_16_sp4_v_b_29_66144),
    .O(seg_17_16_local_g3_5_70017)
  );
  Span4Mux_v4 t2714 (
    .I(seg_17_14_sp4_v_b_5_65652),
    .O(seg_17_16_sp4_v_b_29_66144)
  );
  Span4Mux_v4 t2715 (
    .I(seg_17_10_sp4_h_l_37_54022),
    .O(seg_17_14_sp4_v_b_5_65652)
  );
  LocalMux t2716 (
    .I(seg_17_19_sp4_v_b_41_66637),
    .O(seg_17_19_local_g3_1_70382)
  );
  Span4Mux_v4 t2717 (
    .I(seg_17_18_sp4_v_b_8_66149),
    .O(seg_17_19_sp4_v_b_41_66637)
  );
  Span4Mux_v4 t2718 (
    .I(seg_17_14_sp4_v_b_0_65649),
    .O(seg_17_18_sp4_v_b_8_66149)
  );
  Span4Mux_v4 t2719 (
    .I(seg_17_10_sp4_h_l_37_54022),
    .O(seg_17_14_sp4_v_b_0_65649)
  );
  CascadeMux t272 (
    .I(net_50519),
    .O(net_50519_cascademuxed)
  );
  LocalMux t2720 (
    .I(seg_17_20_sp4_v_b_28_66637),
    .O(seg_17_20_local_g3_4_70508)
  );
  Span4Mux_v4 t2721 (
    .I(seg_17_18_sp4_v_b_8_66149),
    .O(seg_17_20_sp4_v_b_28_66637)
  );
  LocalMux t2722 (
    .I(seg_14_14_sp4_r_v_b_2_57990),
    .O(seg_14_14_local_g1_2_58260)
  );
  Span4Mux_v4 t2723 (
    .I(seg_15_10_sp4_h_r_8_61692),
    .O(seg_14_14_sp4_r_v_b_2_57990)
  );
  LocalMux t2724 (
    .I(seg_14_18_sp4_r_v_b_10_58490),
    .O(seg_14_18_local_g2_2_58760)
  );
  Span4Mux_v4 t2725 (
    .I(seg_15_14_sp4_v_b_2_57990),
    .O(seg_14_18_sp4_r_v_b_10_58490)
  );
  Span4Mux_v4 t2726 (
    .I(seg_15_10_sp4_h_r_8_61692),
    .O(seg_15_14_sp4_v_b_2_57990)
  );
  LocalMux t2727 (
    .I(seg_15_14_sp4_v_b_2_57990),
    .O(seg_15_14_local_g1_2_62090)
  );
  LocalMux t2728 (
    .I(seg_15_18_sp4_v_b_10_58490),
    .O(seg_15_18_local_g0_2_62574)
  );
  Span4Mux_v4 t2729 (
    .I(seg_15_14_sp4_v_b_2_57990),
    .O(seg_15_18_sp4_v_b_10_58490)
  );
  CascadeMux t273 (
    .I(net_50525),
    .O(net_50525_cascademuxed)
  );
  LocalMux t2730 (
    .I(seg_12_19_sp4_v_b_31_47362),
    .O(seg_12_19_local_g3_7_51235)
  );
  Span4Mux_v4 t2731 (
    .I(seg_12_17_sp4_h_r_7_51061),
    .O(seg_12_19_sp4_v_b_31_47362)
  );
  Span4Mux_h4 t2732 (
    .I(seg_16_17_sp4_v_b_7_62192),
    .O(seg_12_17_sp4_h_r_7_51061)
  );
  Span4Mux_v4 t2733 (
    .I(seg_16_13_sp4_v_b_4_61699),
    .O(seg_16_17_sp4_v_b_7_62192)
  );
  LocalMux t2734 (
    .I(seg_15_13_sp4_r_v_b_4_61699),
    .O(seg_15_13_local_g1_4_61969)
  );
  LocalMux t2735 (
    .I(seg_15_15_sp4_r_v_b_31_62192),
    .O(seg_15_15_local_g1_7_62218)
  );
  Span4Mux_v4 t2736 (
    .I(seg_16_13_sp4_v_b_4_61699),
    .O(seg_15_15_sp4_r_v_b_31_62192)
  );
  LocalMux t2737 (
    .I(seg_16_12_sp4_v_b_17_61699),
    .O(seg_16_12_local_g1_1_65674)
  );
  LocalMux t2738 (
    .I(seg_16_13_sp4_v_b_4_61699),
    .O(seg_16_13_local_g0_4_65792)
  );
  LocalMux t2739 (
    .I(seg_16_15_sp4_v_b_31_62192),
    .O(seg_16_15_local_g2_7_66057)
  );
  CascadeMux t274 (
    .I(net_50531),
    .O(net_50531_cascademuxed)
  );
  Span4Mux_v4 t2740 (
    .I(seg_16_13_sp4_v_b_4_61699),
    .O(seg_16_15_sp4_v_b_31_62192)
  );
  LocalMux t2741 (
    .I(seg_16_20_sp4_v_b_23_62689),
    .O(seg_16_20_local_g1_7_66664)
  );
  Span4Mux_v4 t2742 (
    .I(seg_16_17_sp4_v_b_7_62192),
    .O(seg_16_20_sp4_v_b_23_62689)
  );
  LocalMux t2743 (
    .I(seg_17_17_sp4_h_r_18_66383),
    .O(seg_17_17_local_g1_2_70121)
  );
  Span4Mux_h4 t2744 (
    .I(seg_16_17_sp4_v_b_7_62192),
    .O(seg_17_17_sp4_h_r_18_66383)
  );
  LocalMux t2745 (
    .I(seg_16_18_sp4_v_b_5_62313),
    .O(seg_16_18_local_g1_5_66416)
  );
  Span4Mux_v4 t2746 (
    .I(seg_16_14_sp4_v_b_9_61825),
    .O(seg_16_18_sp4_v_b_5_62313)
  );
  Span4Mux_v4 t2747 (
    .I(seg_16_10_sp4_v_b_9_61333),
    .O(seg_16_14_sp4_v_b_9_61825)
  );
  LocalMux t2748 (
    .I(seg_17_14_sp4_h_r_20_66016),
    .O(seg_17_14_local_g1_4_69754)
  );
  Span4Mux_h4 t2749 (
    .I(seg_16_14_sp4_v_b_9_61825),
    .O(seg_17_14_sp4_h_r_20_66016)
  );
  CascadeMux t275 (
    .I(net_50537),
    .O(net_50537_cascademuxed)
  );
  LocalMux t2750 (
    .I(seg_14_12_sp4_r_v_b_0_57742),
    .O(seg_14_12_local_g1_0_58012)
  );
  LocalMux t2751 (
    .I(seg_14_20_sp4_r_v_b_6_58732),
    .O(seg_14_20_local_g1_6_59002)
  );
  Span4Mux_v4 t2752 (
    .I(seg_15_16_sp4_v_b_3_58235),
    .O(seg_14_20_sp4_r_v_b_6_58732)
  );
  Span4Mux_v4 t2753 (
    .I(seg_15_12_sp4_v_b_0_57742),
    .O(seg_15_16_sp4_v_b_3_58235)
  );
  LocalMux t2754 (
    .I(seg_15_15_sp4_v_b_14_58235),
    .O(seg_15_15_local_g0_6_62209)
  );
  Span4Mux_v4 t2755 (
    .I(seg_15_12_sp4_v_b_0_57742),
    .O(seg_15_15_sp4_v_b_14_58235)
  );
  LocalMux t2756 (
    .I(seg_14_13_sp4_r_v_b_5_57868),
    .O(seg_14_13_local_g1_5_58140)
  );
  LocalMux t2757 (
    .I(seg_15_9_sp4_v_b_3_57374),
    .O(seg_15_9_local_g1_3_61476)
  );
  Span4Mux_v4 t2758 (
    .I(seg_15_9_sp4_v_t_42_57870),
    .O(seg_15_9_sp4_v_b_3_57374)
  );
  LocalMux t2759 (
    .I(seg_14_12_neigh_op_bnr_1_57841),
    .O(seg_14_12_local_g1_1_58013)
  );
  CascadeMux t276 (
    .I(net_50543),
    .O(net_50543_cascademuxed)
  );
  LocalMux t2760 (
    .I(seg_14_12_neigh_op_bnr_2_57842),
    .O(seg_14_12_local_g1_2_58014)
  );
  LocalMux t2761 (
    .I(seg_16_12_neigh_op_bnl_4_57844),
    .O(seg_16_12_local_g3_4_65693)
  );
  LocalMux t2762 (
    .I(seg_16_12_neigh_op_bnl_6_57846),
    .O(seg_16_12_local_g2_6_65687)
  );
  LocalMux t2763 (
    .I(seg_14_12_neigh_op_bnr_7_57847),
    .O(seg_14_12_local_g1_7_58019)
  );
  LocalMux t2764 (
    .I(seg_13_13_sp4_r_v_b_29_54284),
    .O(seg_13_13_local_g1_5_54310)
  );
  Span4Mux_v4 t2765 (
    .I(seg_14_11_sp4_h_r_11_57978),
    .O(seg_13_13_sp4_r_v_b_29_54284)
  );
  LocalMux t2766 (
    .I(seg_15_13_sp4_r_v_b_3_61696),
    .O(seg_15_13_local_g1_3_61968)
  );
  LocalMux t2767 (
    .I(seg_15_13_neigh_op_bot_0_57963),
    .O(seg_15_13_local_g0_0_61957)
  );
  LocalMux t2768 (
    .I(seg_14_13_neigh_op_bnr_1_57964),
    .O(seg_14_13_local_g0_1_58128)
  );
  LocalMux t2769 (
    .I(seg_15_13_neigh_op_bot_2_57965),
    .O(seg_15_13_local_g1_2_61967)
  );
  CascadeMux t277 (
    .I(net_50624),
    .O(net_50624_cascademuxed)
  );
  LocalMux t2770 (
    .I(seg_16_13_neigh_op_bnl_3_57966),
    .O(seg_16_13_local_g2_3_65807)
  );
  LocalMux t2771 (
    .I(seg_15_13_neigh_op_bot_4_57967),
    .O(seg_15_13_local_g0_4_61961)
  );
  LocalMux t2772 (
    .I(seg_15_13_neigh_op_bot_5_57968),
    .O(seg_15_13_local_g1_5_61970)
  );
  LocalMux t2773 (
    .I(seg_14_13_neigh_op_bnr_6_57969),
    .O(seg_14_13_local_g1_6_58141)
  );
  LocalMux t2774 (
    .I(seg_14_13_neigh_op_bnr_7_57970),
    .O(seg_14_13_local_g0_7_58134)
  );
  LocalMux t2775 (
    .I(seg_15_12_neigh_op_top_3_58089),
    .O(seg_15_12_local_g0_3_61837)
  );
  LocalMux t2776 (
    .I(seg_15_12_neigh_op_top_4_58090),
    .O(seg_15_12_local_g0_4_61838)
  );
  LocalMux t2777 (
    .I(seg_15_13_lutff_7_out_58093),
    .O(seg_15_13_local_g1_7_61972)
  );
  LocalMux t2778 (
    .I(seg_18_12_sp4_r_v_b_19_73194),
    .O(seg_18_12_local_g3_3_73354)
  );
  Span4Mux_v4 t2779 (
    .I(seg_19_13_sp4_h_l_37_62051),
    .O(seg_18_12_sp4_r_v_b_19_73194)
  );
  CascadeMux t278 (
    .I(net_50636),
    .O(net_50636_cascademuxed)
  );
  LocalMux t2780 (
    .I(seg_19_13_sp4_h_r_8_77111),
    .O(seg_19_13_local_g0_0_77027)
  );
  Span4Mux_h4 t2781 (
    .I(seg_19_13_sp4_h_l_37_62051),
    .O(seg_19_13_sp4_h_r_8_77111)
  );
  LocalMux t2782 (
    .I(seg_18_13_sp4_h_r_47_62053),
    .O(seg_18_13_local_g3_7_73481)
  );
  LocalMux t2783 (
    .I(seg_19_14_sp4_v_b_47_73690),
    .O(seg_19_14_local_g2_7_77152)
  );
  Span4Mux_v4 t2784 (
    .I(seg_19_13_sp4_h_l_47_62053),
    .O(seg_19_14_sp4_v_b_47_73690)
  );
  LocalMux t2785 (
    .I(seg_19_13_sp4_h_r_20_73555),
    .O(seg_19_13_local_g0_4_77031)
  );
  Span4Mux_h4 t2786 (
    .I(seg_18_13_sp4_h_l_36_58222),
    .O(seg_19_13_sp4_h_r_20_73555)
  );
  LocalMux t2787 (
    .I(seg_19_13_sp4_h_r_14_73549),
    .O(seg_19_13_local_g0_6_77033)
  );
  Span4Mux_h4 t2788 (
    .I(seg_18_13_sp4_h_l_42_58230),
    .O(seg_19_13_sp4_h_r_14_73549)
  );
  LocalMux t2789 (
    .I(seg_18_13_sp4_h_r_41_62057),
    .O(seg_18_13_local_g2_1_73467)
  );
  CascadeMux t279 (
    .I(net_50654),
    .O(net_50654_cascademuxed)
  );
  LocalMux t2790 (
    .I(seg_19_13_sp4_h_r_4_77107),
    .O(seg_19_13_local_g1_4_77039)
  );
  Span4Mux_h4 t2791 (
    .I(seg_19_13_sp4_h_l_41_62057),
    .O(seg_19_13_sp4_h_r_4_77107)
  );
  LocalMux t2792 (
    .I(seg_17_14_sp4_h_r_13_66005),
    .O(seg_17_14_local_g0_5_69747)
  );
  Span4Mux_h4 t2793 (
    .I(seg_16_14_sp4_v_b_0_61818),
    .O(seg_17_14_sp4_h_r_13_66005)
  );
  LocalMux t2794 (
    .I(seg_20_14_sp4_h_r_6_80706),
    .O(seg_20_14_local_g1_6_80618)
  );
  Span4Mux_h4 t2795 (
    .I(seg_20_14_sp4_h_l_43_66013),
    .O(seg_20_14_sp4_h_r_6_80706)
  );
  Span4Mux_h4 t2796 (
    .I(seg_16_14_sp4_v_b_6_61824),
    .O(seg_20_14_sp4_h_l_43_66013)
  );
  LocalMux t2797 (
    .I(seg_15_13_neigh_op_top_0_58209),
    .O(seg_15_13_local_g1_0_61965)
  );
  LocalMux t2798 (
    .I(seg_15_14_lutff_0_out_58209),
    .O(seg_15_14_local_g2_0_62096)
  );
  LocalMux t2799 (
    .I(seg_15_13_neigh_op_top_5_58214),
    .O(seg_15_13_local_g0_5_61962)
  );
  CascadeMux t28 (
    .I(net_17421),
    .O(net_17421_cascademuxed)
  );
  CascadeMux t280 (
    .I(net_50666),
    .O(net_50666_cascademuxed)
  );
  LocalMux t2800 (
    .I(seg_15_14_lutff_5_out_58214),
    .O(seg_15_14_local_g2_5_62101)
  );
  LocalMux t2801 (
    .I(seg_20_14_sp4_h_r_27_73672),
    .O(seg_20_14_local_g3_3_80631)
  );
  Span4Mux_h4 t2802 (
    .I(seg_18_14_sp4_h_l_38_58349),
    .O(seg_20_14_sp4_h_r_27_73672)
  );
  LocalMux t2803 (
    .I(seg_17_14_sp4_h_r_26_62178),
    .O(seg_17_14_local_g2_2_69760)
  );
  LocalMux t2804 (
    .I(seg_19_14_sp4_h_r_8_77213),
    .O(seg_19_14_local_g0_0_77129)
  );
  Span4Mux_h4 t2805 (
    .I(seg_19_14_sp4_h_l_45_62184),
    .O(seg_19_14_sp4_h_r_8_77213)
  );
  LocalMux t2806 (
    .I(seg_22_13_sp4_r_v_b_15_88006),
    .O(seg_22_13_local_g2_7_88166)
  );
  Span4Mux_v4 t2807 (
    .I(seg_23_14_sp4_h_l_45_77213),
    .O(seg_22_13_sp4_r_v_b_15_88006)
  );
  Span4Mux_h4 t2808 (
    .I(seg_19_14_sp4_h_l_45_62184),
    .O(seg_23_14_sp4_h_l_45_77213)
  );
  LocalMux t2809 (
    .I(seg_19_15_sp4_h_r_39_66132),
    .O(seg_19_15_local_g2_7_77254)
  );
  CascadeMux t281 (
    .I(net_50759),
    .O(net_50759_cascademuxed)
  );
  Span4Mux_h4 t2810 (
    .I(seg_16_15_sp4_v_b_2_61943),
    .O(seg_19_15_sp4_h_r_39_66132)
  );
  LocalMux t2811 (
    .I(seg_19_15_sp4_h_r_43_66136),
    .O(seg_19_15_local_g3_3_77258)
  );
  Span4Mux_h4 t2812 (
    .I(seg_16_15_sp4_v_b_6_61947),
    .O(seg_19_15_sp4_h_r_43_66136)
  );
  LocalMux t2813 (
    .I(seg_15_12_sp4_r_v_b_31_61823),
    .O(seg_15_12_local_g0_7_61841)
  );
  LocalMux t2814 (
    .I(seg_15_12_sp4_v_b_36_58110),
    .O(seg_15_12_local_g3_4_61862)
  );
  LocalMux t2815 (
    .I(seg_15_12_sp4_v_b_28_57992),
    .O(seg_15_12_local_g2_4_61854)
  );
  LocalMux t2816 (
    .I(seg_15_15_lutff_0_out_58332),
    .O(seg_15_15_local_g3_0_62227)
  );
  LocalMux t2817 (
    .I(seg_15_14_neigh_op_top_1_58333),
    .O(seg_15_14_local_g1_1_62089)
  );
  LocalMux t2818 (
    .I(seg_15_15_lutff_1_out_58333),
    .O(seg_15_15_local_g0_1_62204)
  );
  LocalMux t2819 (
    .I(seg_15_15_lutff_5_out_58337),
    .O(seg_15_15_local_g3_5_62232)
  );
  CascadeMux t282 (
    .I(net_50771),
    .O(net_50771_cascademuxed)
  );
  LocalMux t2820 (
    .I(seg_15_14_neigh_op_top_7_58339),
    .O(seg_15_14_local_g1_7_62095)
  );
  LocalMux t2821 (
    .I(seg_16_15_neigh_op_lft_7_58339),
    .O(seg_16_15_local_g0_7_66041)
  );
  LocalMux t2822 (
    .I(seg_18_15_sp4_h_r_41_62303),
    .O(seg_18_15_local_g2_1_73713)
  );
  LocalMux t2823 (
    .I(seg_19_15_sp4_h_r_0_77305),
    .O(seg_19_15_local_g0_0_77231)
  );
  Span4Mux_h4 t2824 (
    .I(seg_19_15_sp4_h_l_41_62303),
    .O(seg_19_15_sp4_h_r_0_77305)
  );
  LocalMux t2825 (
    .I(seg_18_15_sp4_h_r_45_62307),
    .O(seg_18_15_local_g2_5_73717)
  );
  LocalMux t2826 (
    .I(seg_19_16_sp4_v_b_45_73934),
    .O(seg_19_16_local_g2_5_77354)
  );
  Span4Mux_v4 t2827 (
    .I(seg_19_15_sp4_h_l_45_62307),
    .O(seg_19_16_sp4_v_b_45_73934)
  );
  LocalMux t2828 (
    .I(seg_15_12_sp4_r_v_b_0_61572),
    .O(seg_15_12_local_g1_0_61842)
  );
  Span4Mux_v4 t2829 (
    .I(seg_16_12_sp4_v_t_37_62064),
    .O(seg_15_12_sp4_r_v_b_0_61572)
  );
  CascadeMux t283 (
    .I(net_50777),
    .O(net_50777_cascademuxed)
  );
  LocalMux t2830 (
    .I(seg_15_11_sp4_v_b_15_57744),
    .O(seg_15_11_local_g1_7_61726)
  );
  Span4Mux_v4 t2831 (
    .I(seg_15_12_sp4_v_t_46_58243),
    .O(seg_15_11_sp4_v_b_15_57744)
  );
  LocalMux t2832 (
    .I(seg_15_16_lutff_6_out_58461),
    .O(seg_15_16_local_g2_6_62348)
  );
  LocalMux t2833 (
    .I(seg_13_16_sp4_h_r_2_54764),
    .O(seg_13_16_local_g0_2_54668)
  );
  LocalMux t2834 (
    .I(seg_15_14_sp4_r_v_b_33_62071),
    .O(seg_15_14_local_g0_2_62082)
  );
  LocalMux t2835 (
    .I(seg_15_13_sp4_v_b_37_58234),
    .O(seg_15_13_local_g2_5_61978)
  );
  LocalMux t2836 (
    .I(seg_15_13_sp4_v_b_6_57871),
    .O(seg_15_13_local_g0_6_61963)
  );
  Span4Mux_v4 t2837 (
    .I(seg_15_13_sp4_v_t_38_58358),
    .O(seg_15_13_sp4_v_b_6_57871)
  );
  LocalMux t2838 (
    .I(seg_15_13_sp4_v_b_43_58240),
    .O(seg_15_13_local_g2_3_61976)
  );
  LocalMux t2839 (
    .I(seg_15_17_lutff_0_out_58578),
    .O(seg_15_17_local_g1_0_62457)
  );
  CascadeMux t284 (
    .I(net_50789),
    .O(net_50789_cascademuxed)
  );
  LocalMux t2840 (
    .I(seg_14_17_neigh_op_rgt_2_58580),
    .O(seg_14_17_local_g3_2_58645)
  );
  LocalMux t2841 (
    .I(seg_15_17_lutff_2_out_58580),
    .O(seg_15_17_local_g2_2_62467)
  );
  LocalMux t2842 (
    .I(seg_14_17_neigh_op_rgt_7_58585),
    .O(seg_14_17_local_g3_7_58650)
  );
  LocalMux t2843 (
    .I(seg_15_17_lutff_7_out_58585),
    .O(seg_15_17_local_g2_7_62472)
  );
  LocalMux t2844 (
    .I(seg_13_17_sp4_h_r_4_54889),
    .O(seg_13_17_local_g0_4_54793)
  );
  LocalMux t2845 (
    .I(seg_15_14_sp4_v_b_47_58367),
    .O(seg_15_14_local_g3_7_62111)
  );
  LocalMux t2846 (
    .I(seg_15_15_sp4_v_b_26_58359),
    .O(seg_15_15_local_g2_2_62221)
  );
  LocalMux t2847 (
    .I(seg_15_14_sp4_h_r_4_62180),
    .O(seg_15_14_local_g1_4_62092)
  );
  Span4Mux_h4 t2848 (
    .I(seg_15_14_sp4_v_t_46_58489),
    .O(seg_15_14_sp4_h_r_4_62180)
  );
  LocalMux t2849 (
    .I(seg_15_18_lutff_1_out_58702),
    .O(seg_15_18_local_g0_1_62573)
  );
  LocalMux t2850 (
    .I(seg_16_18_neigh_op_lft_2_58703),
    .O(seg_16_18_local_g0_2_66405)
  );
  LocalMux t2851 (
    .I(seg_15_18_lutff_4_out_58705),
    .O(seg_15_18_local_g3_4_62600)
  );
  LocalMux t2852 (
    .I(seg_15_18_lutff_7_out_58708),
    .O(seg_15_18_local_g0_7_62579)
  );
  LocalMux t2853 (
    .I(seg_18_17_sp4_r_v_b_19_73809),
    .O(seg_18_17_local_g3_3_73969)
  );
  Span4Mux_v4 t2854 (
    .I(seg_19_18_sp4_h_l_37_62666),
    .O(seg_18_17_sp4_r_v_b_19_73809)
  );
  LocalMux t2855 (
    .I(seg_19_18_sp4_h_r_0_77611),
    .O(seg_19_18_local_g1_0_77545)
  );
  Span4Mux_h4 t2856 (
    .I(seg_19_18_sp4_h_l_37_62666),
    .O(seg_19_18_sp4_h_r_0_77611)
  );
  LocalMux t2857 (
    .I(seg_17_18_sp4_h_r_36_58837),
    .O(seg_17_18_local_g2_4_70254)
  );
  LocalMux t2858 (
    .I(seg_19_18_sp4_h_r_12_74160),
    .O(seg_19_18_local_g0_4_77541)
  );
  Span4Mux_h4 t2859 (
    .I(seg_18_18_sp4_h_l_36_58837),
    .O(seg_19_18_sp4_h_r_12_74160)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t286 (
    .carryinitin(),
    .carryinitout(t285)
  );
  LocalMux t2860 (
    .I(seg_15_18_neigh_op_top_0_58824),
    .O(seg_15_18_local_g0_0_62572)
  );
  LocalMux t2861 (
    .I(seg_14_18_neigh_op_tnr_3_58827),
    .O(seg_14_18_local_g2_3_58761)
  );
  LocalMux t2862 (
    .I(seg_14_19_neigh_op_rgt_3_58827),
    .O(seg_14_19_local_g3_3_58892)
  );
  LocalMux t2863 (
    .I(seg_14_20_neigh_op_bnr_3_58827),
    .O(seg_14_20_local_g0_3_58991)
  );
  LocalMux t2864 (
    .I(seg_15_19_lutff_3_out_58827),
    .O(seg_15_19_local_g3_3_62722)
  );
  LocalMux t2865 (
    .I(seg_15_20_neigh_op_bot_3_58827),
    .O(seg_15_20_local_g0_3_62821)
  );
  LocalMux t2866 (
    .I(seg_16_18_neigh_op_tnl_3_58827),
    .O(seg_16_18_local_g3_3_66430)
  );
  LocalMux t2867 (
    .I(seg_15_19_lutff_5_out_58829),
    .O(seg_15_19_local_g3_5_62724)
  );
  LocalMux t2868 (
    .I(seg_15_18_neigh_op_top_6_58830),
    .O(seg_15_18_local_g0_6_62578)
  );
  LocalMux t2869 (
    .I(seg_13_14_sp4_r_v_b_18_54286),
    .O(seg_13_14_local_g3_2_54446)
  );
  CascadeMux t287 (
    .I(net_50876),
    .O(net_50876_cascademuxed)
  );
  Span4Mux_v4 t2870 (
    .I(seg_14_15_sp4_v_t_46_54782),
    .O(seg_13_14_sp4_r_v_b_18_54286)
  );
  Span4Mux_v4 t2871 (
    .I(seg_14_19_sp4_h_r_11_58962),
    .O(seg_14_15_sp4_v_t_46_54782)
  );
  LocalMux t2872 (
    .I(seg_17_17_sp4_r_v_b_29_70098),
    .O(seg_17_17_local_g1_5_70124)
  );
  Span4Mux_v4 t2873 (
    .I(seg_18_19_sp4_h_l_46_58962),
    .O(seg_17_17_sp4_r_v_b_29_70098)
  );
  LocalMux t2874 (
    .I(seg_12_19_sp4_h_r_3_51303),
    .O(seg_12_19_local_g1_3_51215)
  );
  LocalMux t2875 (
    .I(seg_17_19_sp4_h_r_30_62797),
    .O(seg_17_19_local_g2_6_70379)
  );
  LocalMux t2876 (
    .I(seg_17_16_sp4_h_r_23_66253),
    .O(seg_17_16_local_g1_7_70003)
  );
  Span4Mux_h4 t2877 (
    .I(seg_16_16_sp4_v_t_47_62566),
    .O(seg_17_16_sp4_h_r_23_66253)
  );
  LocalMux t2878 (
    .I(seg_17_20_sp4_h_r_17_66749),
    .O(seg_17_20_local_g1_1_70489)
  );
  Span4Mux_h4 t2879 (
    .I(seg_16_20_sp4_v_b_10_62566),
    .O(seg_17_20_sp4_h_r_17_66749)
  );
  CascadeMux t288 (
    .I(net_50906),
    .O(net_50906_cascademuxed)
  );
  LocalMux t2880 (
    .I(seg_16_13_sp4_v_b_34_61951),
    .O(seg_16_13_local_g3_2_65814)
  );
  Span4Mux_v4 t2881 (
    .I(seg_16_15_sp4_v_t_42_62438),
    .O(seg_16_13_sp4_v_b_34_61951)
  );
  LocalMux t2882 (
    .I(seg_16_14_sp4_v_b_23_61951),
    .O(seg_16_14_local_g0_7_65918)
  );
  Span4Mux_v4 t2883 (
    .I(seg_16_15_sp4_v_t_42_62438),
    .O(seg_16_14_sp4_v_b_23_61951)
  );
  LocalMux t2884 (
    .I(seg_16_15_sp4_h_r_0_66128),
    .O(seg_16_15_local_g1_0_66042)
  );
  Span4Mux_h4 t2885 (
    .I(seg_16_15_sp4_v_t_42_62438),
    .O(seg_16_15_sp4_h_r_0_66128)
  );
  LocalMux t2886 (
    .I(seg_17_15_sp4_h_r_18_66137),
    .O(seg_17_15_local_g0_2_69867)
  );
  Span4Mux_h4 t2887 (
    .I(seg_16_15_sp4_v_t_42_62438),
    .O(seg_17_15_sp4_h_r_18_66137)
  );
  LocalMux t2888 (
    .I(seg_12_16_sp4_h_r_16_47105),
    .O(seg_12_16_local_g0_0_50835)
  );
  Span4Mux_h4 t2889 (
    .I(seg_15_16_sp4_v_t_46_58735),
    .O(seg_12_16_sp4_h_r_16_47105)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t289 (
    .carryinitin(net_54740),
    .carryinitout(net_54784)
  );
  LocalMux t2890 (
    .I(seg_13_15_sp4_h_r_24_46975),
    .O(seg_13_15_local_g2_0_54559)
  );
  Span4Mux_h4 t2891 (
    .I(seg_15_15_sp4_v_t_43_58609),
    .O(seg_13_15_sp4_h_r_24_46975)
  );
  LocalMux t2892 (
    .I(seg_14_13_sp4_r_v_b_26_58113),
    .O(seg_14_13_local_g0_2_58129)
  );
  Span4Mux_v4 t2893 (
    .I(seg_15_15_sp4_v_t_43_58609),
    .O(seg_14_13_sp4_r_v_b_26_58113)
  );
  LocalMux t2894 (
    .I(seg_14_13_sp4_r_v_b_30_58117),
    .O(seg_14_13_local_g0_6_58133)
  );
  Span4Mux_v4 t2895 (
    .I(seg_15_15_sp4_v_t_43_58609),
    .O(seg_14_13_sp4_r_v_b_30_58117)
  );
  LocalMux t2896 (
    .I(seg_14_14_sp4_r_v_b_19_58117),
    .O(seg_14_14_local_g3_3_58277)
  );
  Span4Mux_v4 t2897 (
    .I(seg_15_15_sp4_v_t_43_58609),
    .O(seg_14_14_sp4_r_v_b_19_58117)
  );
  LocalMux t2898 (
    .I(seg_14_15_sp4_r_v_b_2_58113),
    .O(seg_14_15_local_g1_2_58383)
  );
  Span4Mux_v4 t2899 (
    .I(seg_15_15_sp4_v_t_43_58609),
    .O(seg_14_15_sp4_r_v_b_2_58113)
  );
  CascadeMux t29 (
    .I(net_17427),
    .O(net_17427_cascademuxed)
  );
  CascadeMux t290 (
    .I(net_50993),
    .O(net_50993_cascademuxed)
  );
  LocalMux t2900 (
    .I(seg_14_16_sp4_r_v_b_43_58609),
    .O(seg_14_16_local_g3_3_58523)
  );
  LocalMux t2901 (
    .I(seg_14_17_sp4_r_v_b_30_58609),
    .O(seg_14_17_local_g1_6_58633)
  );
  LocalMux t2902 (
    .I(seg_15_13_sp4_v_b_26_58113),
    .O(seg_15_13_local_g3_2_61983)
  );
  Span4Mux_v4 t2903 (
    .I(seg_15_15_sp4_v_t_43_58609),
    .O(seg_15_13_sp4_v_b_26_58113)
  );
  LocalMux t2904 (
    .I(seg_15_15_sp4_h_r_11_62300),
    .O(seg_15_15_local_g0_3_62206)
  );
  Span4Mux_h4 t2905 (
    .I(seg_15_15_sp4_v_t_43_58609),
    .O(seg_15_15_sp4_h_r_11_62300)
  );
  LocalMux t2906 (
    .I(seg_15_16_sp4_v_b_43_58609),
    .O(seg_15_16_local_g3_3_62353)
  );
  LocalMux t2907 (
    .I(seg_15_17_sp4_v_b_30_58609),
    .O(seg_15_17_local_g2_6_62471)
  );
  LocalMux t2908 (
    .I(seg_15_19_neigh_op_top_0_58947),
    .O(seg_15_19_local_g1_0_62703)
  );
  LocalMux t2909 (
    .I(seg_15_20_lutff_2_out_58949),
    .O(seg_15_20_local_g1_2_62828)
  );
  CascadeMux t291 (
    .I(net_50999),
    .O(net_50999_cascademuxed)
  );
  LocalMux t2910 (
    .I(seg_14_10_sp4_r_v_b_10_57506),
    .O(seg_14_10_local_g2_2_57776)
  );
  Sp12to4 t2911 (
    .I(seg_15_9_sp12_v_b_23_61435),
    .O(seg_14_10_sp4_r_v_b_10_57506)
  );
  LocalMux t2912 (
    .I(seg_15_10_sp12_v_b_20_61435),
    .O(seg_15_10_local_g3_4_61616)
  );
  LocalMux t2913 (
    .I(seg_13_16_sp4_h_r_11_54763),
    .O(seg_13_16_local_g1_3_54677)
  );
  Span4Mux_h4 t2914 (
    .I(seg_13_16_sp4_v_t_46_51074),
    .O(seg_13_16_sp4_h_r_11_54763)
  );
  Span4Mux_v4 t2915 (
    .I(seg_13_20_sp4_h_r_6_55260),
    .O(seg_13_16_sp4_v_t_46_51074)
  );
  LocalMux t2916 (
    .I(seg_15_20_sp4_r_v_b_3_62557),
    .O(seg_15_20_local_g1_3_62829)
  );
  Span4Mux_v4 t2917 (
    .I(seg_16_20_sp4_h_l_44_51432),
    .O(seg_15_20_sp4_r_v_b_3_62557)
  );
  LocalMux t2918 (
    .I(seg_14_16_sp4_h_r_25_50930),
    .O(seg_14_16_local_g3_1_58521)
  );
  Span4Mux_h4 t2919 (
    .I(seg_16_16_sp4_v_t_36_62555),
    .O(seg_14_16_sp4_h_r_25_50930)
  );
  CascadeMux t292 (
    .I(net_51116),
    .O(net_51116_cascademuxed)
  );
  LocalMux t2920 (
    .I(seg_15_16_sp4_h_r_5_62427),
    .O(seg_15_16_local_g0_5_62331)
  );
  Span4Mux_h4 t2921 (
    .I(seg_15_16_sp4_v_t_37_58726),
    .O(seg_15_16_sp4_h_r_5_62427)
  );
  LocalMux t2922 (
    .I(seg_15_17_sp4_v_b_37_58726),
    .O(seg_15_17_local_g3_5_62478)
  );
  LocalMux t2923 (
    .I(seg_15_18_sp4_v_b_24_58726),
    .O(seg_15_18_local_g2_0_62588)
  );
  LocalMux t2924 (
    .I(seg_13_17_sp4_h_r_27_47226),
    .O(seg_13_17_local_g3_3_54816)
  );
  Span4Mux_h4 t2925 (
    .I(seg_15_17_sp4_v_t_38_58850),
    .O(seg_13_17_sp4_h_r_27_47226)
  );
  LocalMux t2926 (
    .I(seg_15_16_sp4_v_b_19_58363),
    .O(seg_15_16_local_g1_3_62337)
  );
  Span4Mux_v4 t2927 (
    .I(seg_15_17_sp4_v_t_38_58850),
    .O(seg_15_16_sp4_v_b_19_58363)
  );
  LocalMux t2928 (
    .I(seg_14_15_sp4_r_v_b_25_58356),
    .O(seg_14_15_local_g1_1_58382)
  );
  Span4Mux_v4 t2929 (
    .I(seg_15_17_sp4_v_t_40_58852),
    .O(seg_14_15_sp4_r_v_b_25_58356)
  );
  CascadeMux t293 (
    .I(net_51128),
    .O(net_51128_cascademuxed)
  );
  LocalMux t2930 (
    .I(seg_14_15_sp4_v_b_26_54529),
    .O(seg_14_15_local_g2_2_58391)
  );
  Span4Mux_v4 t2931 (
    .I(seg_14_17_sp4_v_t_43_55025),
    .O(seg_14_15_sp4_v_b_26_54529)
  );
  Span4Mux_v4 t2932 (
    .I(seg_14_21_sp4_h_r_1_59206),
    .O(seg_14_17_sp4_v_t_43_55025)
  );
  LocalMux t2933 (
    .I(seg_14_17_sp4_h_r_11_58716),
    .O(seg_14_17_local_g1_3_58630)
  );
  Span4Mux_h4 t2934 (
    .I(seg_14_17_sp4_v_t_43_55025),
    .O(seg_14_17_sp4_h_r_11_58716)
  );
  LocalMux t2935 (
    .I(seg_14_18_sp4_v_b_43_55025),
    .O(seg_14_18_local_g3_3_58769)
  );
  Span4Mux_v4 t2936 (
    .I(seg_14_21_sp4_h_r_1_59206),
    .O(seg_14_18_sp4_v_b_43_55025)
  );
  LocalMux t2937 (
    .I(seg_14_20_sp4_v_b_19_55025),
    .O(seg_14_20_local_g1_3_58999)
  );
  Span4Mux_v4 t2938 (
    .I(seg_14_21_sp4_h_r_1_59206),
    .O(seg_14_20_sp4_v_b_19_55025)
  );
  LocalMux t2939 (
    .I(seg_15_17_sp4_h_r_19_58721),
    .O(seg_15_17_local_g1_3_62460)
  );
  CascadeMux t294 (
    .I(net_51251),
    .O(net_51251_cascademuxed)
  );
  Span4Mux_h4 t2940 (
    .I(seg_14_17_sp4_v_t_43_55025),
    .O(seg_15_17_sp4_h_r_19_58721)
  );
  LocalMux t2941 (
    .I(seg_17_19_sp4_v_b_34_66520),
    .O(seg_17_19_local_g2_2_70375)
  );
  Span4Mux_v4 t2942 (
    .I(seg_17_21_sp4_h_l_41_55381),
    .O(seg_17_19_sp4_v_b_34_66520)
  );
  LocalMux t2943 (
    .I(seg_17_21_sp4_v_b_10_66520),
    .O(seg_17_21_local_g0_2_70605)
  );
  Span4Mux_v4 t2944 (
    .I(seg_17_21_sp4_h_l_41_55381),
    .O(seg_17_21_sp4_v_b_10_66520)
  );
  LocalMux t2945 (
    .I(seg_12_17_sp4_h_r_2_51056),
    .O(seg_12_17_local_g0_2_50960)
  );
  Span4Mux_h4 t2946 (
    .I(seg_12_17_sp4_v_t_44_47364),
    .O(seg_12_17_sp4_h_r_2_51056)
  );
  Span4Mux_v4 t2947 (
    .I(seg_12_21_sp4_h_r_9_51555),
    .O(seg_12_17_sp4_v_t_44_47364)
  );
  LocalMux t2948 (
    .I(seg_12_19_sp4_v_b_26_47359),
    .O(seg_12_19_local_g2_2_51222)
  );
  Span4Mux_v4 t2949 (
    .I(seg_12_21_sp4_h_r_9_51555),
    .O(seg_12_19_sp4_v_b_26_47359)
  );
  CascadeMux t295 (
    .I(net_51263),
    .O(net_51263_cascademuxed)
  );
  LocalMux t2950 (
    .I(seg_15_19_sp4_r_v_b_27_62680),
    .O(seg_15_19_local_g1_3_62706)
  );
  Span4Mux_v4 t2951 (
    .I(seg_16_21_sp4_h_l_44_51555),
    .O(seg_15_19_sp4_r_v_b_27_62680)
  );
  LocalMux t2952 (
    .I(seg_12_16_sp4_v_b_35_46997),
    .O(seg_12_16_local_g3_3_50862)
  );
  Span4Mux_v4 t2953 (
    .I(seg_12_18_sp4_h_r_6_51183),
    .O(seg_12_16_sp4_v_b_35_46997)
  );
  Span4Mux_h4 t2954 (
    .I(seg_16_18_sp4_v_t_37_62802),
    .O(seg_12_18_sp4_h_r_6_51183)
  );
  LocalMux t2955 (
    .I(seg_16_16_sp4_v_b_27_62311),
    .O(seg_16_16_local_g3_3_66184)
  );
  Span4Mux_v4 t2956 (
    .I(seg_16_18_sp4_v_t_37_62802),
    .O(seg_16_16_sp4_v_b_27_62311)
  );
  LocalMux t2957 (
    .I(seg_14_16_sp4_r_v_b_33_58487),
    .O(seg_14_16_local_g0_2_58498)
  );
  Span4Mux_v4 t2958 (
    .I(seg_15_18_sp4_v_t_36_58971),
    .O(seg_14_16_sp4_r_v_b_33_58487)
  );
  LocalMux t2959 (
    .I(seg_16_18_sp4_h_r_19_62674),
    .O(seg_16_18_local_g1_3_66414)
  );
  CascadeMux t296 (
    .I(net_51485),
    .O(net_51485_cascademuxed)
  );
  Span4Mux_h4 t2960 (
    .I(seg_15_18_sp4_v_t_36_58971),
    .O(seg_16_18_sp4_h_r_19_62674)
  );
  LocalMux t2961 (
    .I(seg_15_22_lutff_4_out_59197),
    .O(seg_15_22_local_g0_4_63068)
  );
  LocalMux t2962 (
    .I(seg_15_23_neigh_op_bot_5_59198),
    .O(seg_15_23_local_g1_5_63200)
  );
  LocalMux t2963 (
    .I(seg_13_16_sp4_h_r_27_47103),
    .O(seg_13_16_local_g2_3_54685)
  );
  Span4Mux_h4 t2964 (
    .I(seg_15_16_sp4_v_t_38_58727),
    .O(seg_13_16_sp4_h_r_27_47103)
  );
  Span4Mux_v4 t2965 (
    .I(seg_15_20_sp4_v_t_37_59218),
    .O(seg_15_16_sp4_v_t_38_58727)
  );
  LocalMux t2966 (
    .I(seg_15_16_sp4_v_b_32_58488),
    .O(seg_15_16_local_g3_0_62350)
  );
  Span4Mux_v4 t2967 (
    .I(seg_15_18_sp4_v_t_45_58980),
    .O(seg_15_16_sp4_v_b_32_58488)
  );
  LocalMux t2968 (
    .I(seg_15_23_lutff_1_out_59317),
    .O(seg_15_23_local_g2_1_63204)
  );
  LocalMux t2969 (
    .I(seg_15_20_sp4_r_v_b_36_62924),
    .O(seg_15_20_local_g2_4_62838)
  );
  CascadeMux t297 (
    .I(net_51521),
    .O(net_51521_cascademuxed)
  );
  Span4Mux_v4 t2970 (
    .I(seg_16_23_sp4_h_l_42_51799),
    .O(seg_15_20_sp4_r_v_b_36_62924)
  );
  LocalMux t2971 (
    .I(seg_15_20_sp4_v_b_47_59105),
    .O(seg_15_20_local_g3_7_62849)
  );
  LocalMux t2972 (
    .I(seg_15_21_sp4_v_b_34_59105),
    .O(seg_15_21_local_g3_2_62967)
  );
  LocalMux t2973 (
    .I(seg_15_20_sp4_h_r_8_62922),
    .O(seg_15_20_local_g0_0_62818)
  );
  Span4Mux_h4 t2974 (
    .I(seg_15_20_sp4_v_t_38_59219),
    .O(seg_15_20_sp4_h_r_8_62922)
  );
  LocalMux t2975 (
    .I(seg_15_20_sp4_r_v_b_18_62684),
    .O(seg_15_20_local_g3_2_62844)
  );
  Span4Mux_v4 t2976 (
    .I(seg_16_21_sp4_v_t_46_63180),
    .O(seg_15_20_sp4_r_v_b_18_62684)
  );
  LocalMux t2977 (
    .I(seg_15_21_sp4_r_v_b_7_62684),
    .O(seg_15_21_local_g1_7_62956)
  );
  Span4Mux_v4 t2978 (
    .I(seg_16_21_sp4_v_t_46_63180),
    .O(seg_15_21_sp4_r_v_b_7_62684)
  );
  LocalMux t2979 (
    .I(seg_15_22_sp4_r_v_b_19_62931),
    .O(seg_15_22_local_g3_3_63091)
  );
  CascadeMux t298 (
    .I(net_51527),
    .O(net_51527_cascademuxed)
  );
  Span4Mux_v4 t2980 (
    .I(seg_16_23_sp4_v_t_38_63418),
    .O(seg_15_22_sp4_r_v_b_19_62931)
  );
  LocalMux t2981 (
    .I(seg_15_23_sp4_v_b_34_59351),
    .O(seg_15_23_local_g2_2_63205)
  );
  LocalMux t2982 (
    .I(seg_15_20_sp4_v_b_40_59098),
    .O(seg_15_20_local_g2_0_62834)
  );
  Span4Mux_v4 t2983 (
    .I(seg_15_23_sp4_v_t_39_59589),
    .O(seg_15_20_sp4_v_b_40_59098)
  );
  LocalMux t2984 (
    .I(seg_14_27_sp4_r_v_b_10_59597),
    .O(seg_14_27_local_g2_2_59867)
  );
  LocalMux t2985 (
    .I(seg_14_28_neigh_op_rgt_0_59931),
    .O(seg_14_28_local_g2_0_59988)
  );
  LocalMux t2986 (
    .I(seg_15_27_neigh_op_top_4_59935),
    .O(seg_15_27_local_g0_4_63683)
  );
  LocalMux t2987 (
    .I(seg_15_28_lutff_5_out_59936),
    .O(seg_15_28_local_g0_5_63807)
  );
  LocalMux t2988 (
    .I(seg_12_27_sp4_r_v_b_19_52055),
    .O(seg_12_27_local_g3_3_52215)
  );
  Span4Mux_v4 t2989 (
    .I(seg_13_28_sp4_h_r_6_56244),
    .O(seg_12_27_sp4_r_v_b_19_52055)
  );
  CascadeMux t299 (
    .I(net_52223),
    .O(net_52223_cascademuxed)
  );
  LocalMux t2990 (
    .I(seg_13_27_sp4_v_b_19_52055),
    .O(seg_13_27_local_g1_3_56030)
  );
  Span4Mux_v4 t2991 (
    .I(seg_13_28_sp4_h_r_6_56244),
    .O(seg_13_27_sp4_v_b_19_52055)
  );
  LocalMux t2992 (
    .I(seg_12_28_sp4_h_r_11_52408),
    .O(seg_12_28_local_g1_3_52322)
  );
  LocalMux t2993 (
    .I(seg_15_25_sp4_v_b_3_59342),
    .O(seg_15_25_local_g1_3_63444)
  );
  Span4Mux_v4 t2994 (
    .I(seg_15_25_sp4_v_t_42_59838),
    .O(seg_15_25_sp4_v_b_3_59342)
  );
  LocalMux t2995 (
    .I(seg_15_29_lutff_5_out_60059),
    .O(seg_15_29_local_g3_5_63954)
  );
  LocalMux t2996 (
    .I(seg_17_31_span4_horz_r_5_68032),
    .O(seg_17_31_local_g1_5_71859)
  );
  IoSpan4Mux t2997 (
    .I(seg_16_31_span4_vert_7_63914),
    .O(seg_17_31_span4_horz_r_5_68032)
  );
  LocalMux t2998 (
    .I(seg_16_2_lutff_1_out_60528),
    .O(seg_16_2_local_g1_1_64444)
  );
  LocalMux t2999 (
    .I(seg_16_2_lutff_2_out_60529),
    .O(seg_16_2_local_g3_2_64461)
  );
  CascadeMux t3 (
    .I(net_12213),
    .O(net_12213_cascademuxed)
  );
  CascadeMux t30 (
    .I(net_17433),
    .O(net_17433_cascademuxed)
  );
  CascadeMux t300 (
    .I(net_52229),
    .O(net_52229_cascademuxed)
  );
  LocalMux t3000 (
    .I(seg_15_3_neigh_op_bnr_5_60532),
    .O(seg_15_3_local_g1_5_60740)
  );
  LocalMux t3001 (
    .I(seg_17_5_neigh_op_lft_2_60934),
    .O(seg_17_5_local_g1_2_68645)
  );
  LocalMux t3002 (
    .I(seg_17_5_neigh_op_lft_3_60935),
    .O(seg_17_5_local_g0_3_68638)
  );
  LocalMux t3003 (
    .I(seg_17_5_neigh_op_lft_4_60936),
    .O(seg_17_5_local_g1_4_68647)
  );
  LocalMux t3004 (
    .I(seg_17_5_neigh_op_lft_5_60937),
    .O(seg_17_5_local_g1_5_68648)
  );
  LocalMux t3005 (
    .I(seg_17_5_neigh_op_lft_6_60938),
    .O(seg_17_5_local_g1_6_68649)
  );
  LocalMux t3006 (
    .I(seg_17_5_neigh_op_lft_7_60939),
    .O(seg_17_5_local_g1_7_68650)
  );
  LocalMux t3007 (
    .I(seg_17_6_neigh_op_lft_0_61055),
    .O(seg_17_6_local_g1_0_68766)
  );
  LocalMux t3008 (
    .I(seg_15_9_neigh_op_rgt_2_61426),
    .O(seg_15_9_local_g2_2_61483)
  );
  LocalMux t3009 (
    .I(seg_16_9_lutff_2_out_61426),
    .O(seg_16_9_local_g0_2_65298)
  );
  CascadeMux t301 (
    .I(net_52241),
    .O(net_52241_cascademuxed)
  );
  LocalMux t3010 (
    .I(seg_16_9_lutff_3_out_61427),
    .O(seg_16_9_local_g2_3_65315)
  );
  LocalMux t3011 (
    .I(seg_16_9_lutff_4_out_61428),
    .O(seg_16_9_local_g1_4_65308)
  );
  LocalMux t3012 (
    .I(seg_15_9_neigh_op_rgt_5_61429),
    .O(seg_15_9_local_g2_5_61486)
  );
  LocalMux t3013 (
    .I(seg_15_10_neigh_op_bnr_6_61430),
    .O(seg_15_10_local_g0_6_61594)
  );
  LocalMux t3014 (
    .I(seg_16_9_lutff_6_out_61430),
    .O(seg_16_9_local_g0_6_65302)
  );
  GlobalMux t3015 (
    .I(seg_6_31_local_g0_7_29714_i3),
    .O(seg_5_20_glb_netwk_3_8)
  );
  gio2CtrlBuf t3016 (
    .I(seg_6_31_local_g0_7_29714_i2),
    .O(seg_6_31_local_g0_7_29714_i3)
  );
  ICE_GB t3017 (
    .GLOBALBUFFEROUTPUT(seg_6_31_local_g0_7_29714_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_6_31_local_g0_7_29714_i1)
  );
  IoInMux t3018 (
    .I(seg_6_31_local_g0_7_29714),
    .O(seg_6_31_local_g0_7_29714_i1)
  );
  LocalMux t3019 (
    .I(seg_6_31_span4_vert_15_26357),
    .O(seg_6_31_local_g0_7_29714)
  );
  CascadeMux t302 (
    .I(net_52352),
    .O(net_52352_cascademuxed)
  );
  Span4Mux_v4 t3020 (
    .I(seg_6_28_sp4_h_r_2_29465),
    .O(seg_6_31_span4_vert_15_26357)
  );
  Sp12to4 t3021 (
    .I(seg_7_28_sp12_h_r_6_22385),
    .O(seg_6_28_sp4_h_r_2_29465)
  );
  Span12Mux_h12 t3022 (
    .I(seg_16_28_sp12_v_b_1_66249),
    .O(seg_7_28_sp12_h_r_6_22385)
  );
  Span12Mux_v12 t3023 (
    .I(seg_16_16_sp12_v_b_1_64773),
    .O(seg_16_28_sp12_v_b_1_66249)
  );
  LocalMux t3024 (
    .I(seg_15_9_sp4_r_v_b_36_61571),
    .O(seg_15_9_local_g2_4_61485)
  );
  LocalMux t3025 (
    .I(seg_15_11_sp4_r_v_b_20_61579),
    .O(seg_15_11_local_g3_4_61739)
  );
  LocalMux t3026 (
    .I(seg_15_10_neigh_op_rgt_5_61552),
    .O(seg_15_10_local_g2_5_61609)
  );
  LocalMux t3027 (
    .I(seg_15_11_neigh_op_bnr_5_61552),
    .O(seg_15_11_local_g1_5_61724)
  );
  LocalMux t3028 (
    .I(seg_15_11_neigh_op_rgt_0_61670),
    .O(seg_15_11_local_g3_0_61735)
  );
  LocalMux t3029 (
    .I(seg_15_11_neigh_op_rgt_1_61671),
    .O(seg_15_11_local_g3_1_61736)
  );
  CascadeMux t303 (
    .I(net_52358),
    .O(net_52358_cascademuxed)
  );
  LocalMux t3030 (
    .I(seg_15_11_neigh_op_rgt_4_61674),
    .O(seg_15_11_local_g2_4_61731)
  );
  LocalMux t3031 (
    .I(seg_16_11_lutff_5_out_61675),
    .O(seg_16_11_local_g0_5_65547)
  );
  LocalMux t3032 (
    .I(seg_16_12_neigh_op_bot_5_61675),
    .O(seg_16_12_local_g1_5_65678)
  );
  LocalMux t3033 (
    .I(seg_16_11_neigh_op_top_2_61795),
    .O(seg_16_11_local_g1_2_65552)
  );
  LocalMux t3034 (
    .I(seg_16_12_lutff_2_out_61795),
    .O(seg_16_12_local_g1_2_65675)
  );
  LocalMux t3035 (
    .I(seg_21_12_sp4_h_r_13_80452),
    .O(seg_21_12_local_g1_5_84202)
  );
  Span4Mux_h4 t3036 (
    .I(seg_20_12_sp4_h_l_37_65759),
    .O(seg_21_12_sp4_h_r_13_80452)
  );
  LocalMux t3037 (
    .I(seg_19_16_sp4_v_b_1_73556),
    .O(seg_19_16_local_g1_1_77342)
  );
  Span4Mux_v4 t3038 (
    .I(seg_19_12_sp4_h_l_36_61929),
    .O(seg_19_16_sp4_v_b_1_73556)
  );
  LocalMux t3039 (
    .I(seg_21_12_sp4_h_r_28_77005),
    .O(seg_21_12_local_g3_4_84217)
  );
  CascadeMux t304 (
    .I(net_53144),
    .O(net_53144_cascademuxed)
  );
  Span4Mux_h4 t3040 (
    .I(seg_19_12_sp4_h_l_36_61929),
    .O(seg_21_12_sp4_h_r_28_77005)
  );
  LocalMux t3041 (
    .I(seg_20_11_sp4_v_b_15_76708),
    .O(seg_20_11_local_g0_7_80242)
  );
  Span4Mux_v4 t3042 (
    .I(seg_20_12_sp4_h_l_39_65763),
    .O(seg_20_11_sp4_v_b_15_76708)
  );
  LocalMux t3043 (
    .I(seg_10_12_sp4_h_r_16_38951),
    .O(seg_10_12_local_g0_0_42681)
  );
  Span4Mux_h4 t3044 (
    .I(seg_13_12_sp4_h_r_5_54275),
    .O(seg_10_12_sp4_h_r_16_38951)
  );
  LocalMux t3045 (
    .I(seg_19_14_sp4_h_r_29_69843),
    .O(seg_19_14_local_g3_5_77158)
  );
  Span4Mux_h4 t3046 (
    .I(seg_17_14_sp4_v_b_11_65658),
    .O(seg_19_14_sp4_h_r_29_69843)
  );
  LocalMux t3047 (
    .I(seg_19_14_sp4_h_r_39_66009),
    .O(seg_19_14_local_g3_7_77160)
  );
  Span4Mux_h4 t3048 (
    .I(seg_16_14_sp4_v_b_8_61826),
    .O(seg_19_14_sp4_h_r_39_66009)
  );
  LocalMux t3049 (
    .I(seg_16_15_sp4_v_b_7_61946),
    .O(seg_16_15_local_g1_7_66049)
  );
  CascadeMux t305 (
    .I(net_53225),
    .O(net_53225_cascademuxed)
  );
  LocalMux t3050 (
    .I(seg_17_13_neigh_op_lft_0_61916),
    .O(seg_17_13_local_g0_0_69619)
  );
  LocalMux t3051 (
    .I(seg_16_13_lutff_2_out_61918),
    .O(seg_16_13_local_g0_2_65790)
  );
  LocalMux t3052 (
    .I(seg_17_13_neigh_op_lft_3_61919),
    .O(seg_17_13_local_g1_3_69630)
  );
  LocalMux t3053 (
    .I(seg_16_12_neigh_op_top_4_61920),
    .O(seg_16_12_local_g1_4_65677)
  );
  LocalMux t3054 (
    .I(seg_19_13_sp4_h_r_41_65888),
    .O(seg_19_13_local_g2_1_77044)
  );
  LocalMux t3055 (
    .I(seg_16_15_neigh_op_bot_1_62040),
    .O(seg_16_15_local_g0_1_66035)
  );
  LocalMux t3056 (
    .I(seg_16_13_neigh_op_top_5_62044),
    .O(seg_16_13_local_g1_5_65801)
  );
  LocalMux t3057 (
    .I(seg_16_14_lutff_7_out_62046),
    .O(seg_16_14_local_g3_7_65942)
  );
  LocalMux t3058 (
    .I(seg_16_12_sp4_v_b_38_61942),
    .O(seg_16_12_local_g3_6_65695)
  );
  LocalMux t3059 (
    .I(seg_16_15_lutff_0_out_62162),
    .O(seg_16_15_local_g2_0_66050)
  );
  CascadeMux t306 (
    .I(net_53231),
    .O(net_53231_cascademuxed)
  );
  LocalMux t3060 (
    .I(seg_16_15_lutff_3_out_62165),
    .O(seg_16_15_local_g3_3_66061)
  );
  LocalMux t3061 (
    .I(seg_16_15_lutff_7_out_62169),
    .O(seg_16_15_local_g3_7_66065)
  );
  LocalMux t3062 (
    .I(seg_18_15_sp4_h_r_34_66130),
    .O(seg_18_15_local_g3_2_73722)
  );
  LocalMux t3063 (
    .I(seg_19_15_sp4_h_r_9_77316),
    .O(seg_19_15_local_g1_1_77240)
  );
  Span4Mux_h4 t3064 (
    .I(seg_19_15_sp4_h_l_36_62298),
    .O(seg_19_15_sp4_h_r_9_77316)
  );
  LocalMux t3065 (
    .I(seg_22_15_sp4_h_r_44_77316),
    .O(seg_22_15_local_g3_4_88417)
  );
  Span4Mux_h4 t3066 (
    .I(seg_19_15_sp4_h_l_36_62298),
    .O(seg_22_15_sp4_h_r_44_77316)
  );
  LocalMux t3067 (
    .I(seg_18_15_sp4_h_r_28_66134),
    .O(seg_18_15_local_g3_4_73724)
  );
  LocalMux t3068 (
    .I(seg_16_11_sp4_r_v_b_16_65406),
    .O(seg_16_11_local_g3_0_65566)
  );
  Span4Mux_v4 t3069 (
    .I(seg_17_12_sp4_v_t_39_65897),
    .O(seg_16_11_sp4_r_v_b_16_65406)
  );
  CascadeMux t307 (
    .I(net_53237),
    .O(net_53237_cascademuxed)
  );
  LocalMux t3070 (
    .I(seg_19_16_sp4_h_r_32_70092),
    .O(seg_19_16_local_g3_0_77357)
  );
  Span4Mux_h4 t3071 (
    .I(seg_17_16_sp4_v_b_8_65903),
    .O(seg_19_16_sp4_h_r_32_70092)
  );
  LocalMux t3072 (
    .I(seg_19_16_sp4_r_v_b_15_77218),
    .O(seg_19_16_local_g2_7_77356)
  );
  Span4Mux_v4 t3073 (
    .I(seg_20_17_sp4_h_l_39_66378),
    .O(seg_19_16_sp4_r_v_b_15_77218)
  );
  Span4Mux_h4 t3074 (
    .I(seg_16_17_sp4_v_b_2_62189),
    .O(seg_20_17_sp4_h_l_39_66378)
  );
  LocalMux t3075 (
    .I(seg_16_12_sp4_v_b_45_61949),
    .O(seg_16_12_local_g2_5_65686)
  );
  LocalMux t3076 (
    .I(seg_17_17_neigh_op_bnl_1_62286),
    .O(seg_17_17_local_g3_1_70136)
  );
  LocalMux t3077 (
    .I(seg_15_16_neigh_op_rgt_2_62287),
    .O(seg_15_16_local_g2_2_62344)
  );
  LocalMux t3078 (
    .I(seg_16_15_neigh_op_top_2_62287),
    .O(seg_16_15_local_g0_2_66036)
  );
  LocalMux t3079 (
    .I(seg_16_19_sp4_v_b_21_62564),
    .O(seg_16_19_local_g0_5_66531)
  );
  CascadeMux t308 (
    .I(net_53255),
    .O(net_53255_cascademuxed)
  );
  Span4Mux_v4 t3080 (
    .I(seg_16_16_sp4_h_r_2_66255),
    .O(seg_16_19_sp4_v_b_21_62564)
  );
  LocalMux t3081 (
    .I(seg_13_13_sp4_h_r_0_54391),
    .O(seg_13_13_local_g0_0_54297)
  );
  Span4Mux_h4 t3082 (
    .I(seg_17_13_sp4_v_t_43_66024),
    .O(seg_13_13_sp4_h_r_0_54391)
  );
  LocalMux t3083 (
    .I(seg_17_12_sp4_v_b_15_65528),
    .O(seg_17_12_local_g0_7_69503)
  );
  Span4Mux_v4 t3084 (
    .I(seg_17_13_sp4_v_t_43_66024),
    .O(seg_17_12_sp4_v_b_15_65528)
  );
  LocalMux t3085 (
    .I(seg_11_10_sp4_r_v_b_26_46252),
    .O(seg_11_10_local_g1_2_46276)
  );
  Span4Mux_v4 t3086 (
    .I(seg_12_12_sp4_h_r_2_50441),
    .O(seg_11_10_sp4_r_v_b_26_46252)
  );
  Span4Mux_h4 t3087 (
    .I(seg_16_12_sp4_v_t_39_62066),
    .O(seg_12_12_sp4_h_r_2_50441)
  );
  LocalMux t3088 (
    .I(seg_13_12_sp4_h_r_15_50441),
    .O(seg_13_12_local_g1_7_54189)
  );
  Span4Mux_h4 t3089 (
    .I(seg_16_12_sp4_v_t_39_62066),
    .O(seg_13_12_sp4_h_r_15_50441)
  );
  CascadeMux t309 (
    .I(net_53267),
    .O(net_53267_cascademuxed)
  );
  LocalMux t3090 (
    .I(seg_16_14_sp4_v_b_26_62066),
    .O(seg_16_14_local_g3_2_65937)
  );
  LocalMux t3091 (
    .I(seg_11_14_sp4_r_v_b_3_46497),
    .O(seg_11_14_local_g1_3_46769)
  );
  Span4Mux_v4 t3092 (
    .I(seg_12_14_sp4_h_r_10_50685),
    .O(seg_11_14_sp4_r_v_b_3_46497)
  );
  Span4Mux_h4 t3093 (
    .I(seg_16_14_sp4_v_t_47_62320),
    .O(seg_12_14_sp4_h_r_10_50685)
  );
  LocalMux t3094 (
    .I(seg_17_17_neigh_op_lft_1_62409),
    .O(seg_17_17_local_g1_1_70120)
  );
  LocalMux t3095 (
    .I(seg_17_18_neigh_op_lft_2_62533),
    .O(seg_17_18_local_g0_2_70236)
  );
  LocalMux t3096 (
    .I(seg_16_18_lutff_3_out_62534),
    .O(seg_16_18_local_g2_3_66422)
  );
  LocalMux t3097 (
    .I(seg_16_18_lutff_4_out_62535),
    .O(seg_16_18_local_g1_4_66415)
  );
  LocalMux t3098 (
    .I(seg_19_18_sp4_h_r_41_66503),
    .O(seg_19_18_local_g3_1_77562)
  );
  LocalMux t3099 (
    .I(seg_17_19_neigh_op_lft_1_62655),
    .O(seg_17_19_local_g0_1_70358)
  );
  CascadeMux t31 (
    .I(net_17514),
    .O(net_17514_cascademuxed)
  );
  CascadeMux t310 (
    .I(net_53735),
    .O(net_53735_cascademuxed)
  );
  LocalMux t3100 (
    .I(seg_16_19_lutff_3_out_62657),
    .O(seg_16_19_local_g1_3_66537)
  );
  LocalMux t3101 (
    .I(seg_16_19_lutff_4_out_62658),
    .O(seg_16_19_local_g3_4_66554)
  );
  LocalMux t3102 (
    .I(seg_16_18_neigh_op_top_5_62659),
    .O(seg_16_18_local_g0_5_66408)
  );
  LocalMux t3103 (
    .I(seg_17_19_neigh_op_lft_6_62660),
    .O(seg_17_19_local_g0_6_70363)
  );
  LocalMux t3104 (
    .I(seg_16_19_lutff_7_out_62661),
    .O(seg_16_19_local_g3_7_66557)
  );
  LocalMux t3105 (
    .I(seg_16_20_lutff_1_out_62778),
    .O(seg_16_20_local_g3_1_66674)
  );
  LocalMux t3106 (
    .I(seg_16_19_neigh_op_top_2_62779),
    .O(seg_16_19_local_g0_2_66528)
  );
  LocalMux t3107 (
    .I(seg_17_19_neigh_op_tnl_3_62780),
    .O(seg_17_19_local_g2_3_70376)
  );
  LocalMux t3108 (
    .I(seg_16_20_lutff_4_out_62781),
    .O(seg_16_20_local_g0_4_66653)
  );
  LocalMux t3109 (
    .I(seg_17_20_neigh_op_lft_5_62782),
    .O(seg_17_20_local_g1_5_70493)
  );
  CascadeMux t311 (
    .I(net_53741),
    .O(net_53741_cascademuxed)
  );
  LocalMux t3110 (
    .I(seg_16_19_neigh_op_top_7_62784),
    .O(seg_16_19_local_g0_7_66533)
  );
  LocalMux t3111 (
    .I(seg_16_20_neigh_op_top_7_62907),
    .O(seg_16_20_local_g0_7_66656)
  );
  LocalMux t3112 (
    .I(seg_15_28_neigh_op_rgt_1_63762),
    .O(seg_15_28_local_g2_1_63819)
  );
  LocalMux t3113 (
    .I(seg_15_29_neigh_op_bnr_1_63762),
    .O(seg_15_29_local_g1_1_63934)
  );
  LocalMux t3114 (
    .I(seg_16_28_lutff_1_out_63762),
    .O(seg_16_28_local_g1_1_67642)
  );
  LocalMux t3115 (
    .I(seg_16_28_lutff_1_out_63762),
    .O(seg_16_28_local_g2_1_67650)
  );
  LocalMux t3116 (
    .I(seg_16_29_neigh_op_bot_1_63762),
    .O(seg_16_29_local_g0_1_67757)
  );
  LocalMux t3117 (
    .I(seg_16_29_neigh_op_bot_1_63762),
    .O(seg_16_29_local_g1_1_67765)
  );
  LocalMux t3118 (
    .I(seg_17_29_neigh_op_bnl_1_63762),
    .O(seg_17_29_local_g2_1_71604)
  );
  LocalMux t3119 (
    .I(seg_16_28_lutff_2_out_63763),
    .O(seg_16_28_local_g1_2_67643)
  );
  CascadeMux t312 (
    .I(net_53747),
    .O(net_53747_cascademuxed)
  );
  LocalMux t3120 (
    .I(seg_15_28_neigh_op_rgt_3_63764),
    .O(seg_15_28_local_g3_3_63829)
  );
  LocalMux t3121 (
    .I(seg_15_29_neigh_op_bnr_3_63764),
    .O(seg_15_29_local_g0_3_63928)
  );
  LocalMux t3122 (
    .I(seg_16_28_lutff_3_out_63764),
    .O(seg_16_28_local_g3_3_67660)
  );
  LocalMux t3123 (
    .I(seg_16_29_neigh_op_bot_3_63764),
    .O(seg_16_29_local_g1_3_67767)
  );
  LocalMux t3124 (
    .I(seg_17_29_neigh_op_bnl_3_63764),
    .O(seg_17_29_local_g3_3_71614)
  );
  LocalMux t3125 (
    .I(seg_15_28_neigh_op_rgt_5_63766),
    .O(seg_15_28_local_g2_5_63823)
  );
  LocalMux t3126 (
    .I(seg_15_28_neigh_op_rgt_5_63766),
    .O(seg_15_28_local_g3_5_63831)
  );
  LocalMux t3127 (
    .I(seg_15_29_neigh_op_bnr_5_63766),
    .O(seg_15_29_local_g0_5_63930)
  );
  LocalMux t3128 (
    .I(seg_15_29_neigh_op_bnr_5_63766),
    .O(seg_15_29_local_g1_5_63938)
  );
  LocalMux t3129 (
    .I(seg_16_28_lutff_5_out_63766),
    .O(seg_16_28_local_g2_5_67654)
  );
  CascadeMux t313 (
    .I(net_53753),
    .O(net_53753_cascademuxed)
  );
  LocalMux t3130 (
    .I(seg_16_29_neigh_op_bot_5_63766),
    .O(seg_16_29_local_g0_5_67761)
  );
  LocalMux t3131 (
    .I(seg_17_29_neigh_op_bnl_5_63766),
    .O(seg_17_29_local_g2_5_71608)
  );
  LocalMux t3132 (
    .I(seg_15_28_neigh_op_rgt_6_63767),
    .O(seg_15_28_local_g2_6_63824)
  );
  LocalMux t3133 (
    .I(seg_15_29_neigh_op_bnr_6_63767),
    .O(seg_15_29_local_g1_6_63939)
  );
  LocalMux t3134 (
    .I(seg_16_28_lutff_6_out_63767),
    .O(seg_16_28_local_g1_6_67647)
  );
  LocalMux t3135 (
    .I(seg_16_29_neigh_op_bot_6_63767),
    .O(seg_16_29_local_g1_6_67770)
  );
  LocalMux t3136 (
    .I(seg_17_29_neigh_op_bnl_6_63767),
    .O(seg_17_29_local_g2_6_71609)
  );
  LocalMux t3137 (
    .I(seg_16_28_lutff_7_out_63768),
    .O(seg_16_28_local_g2_7_67656)
  );
  LocalMux t3138 (
    .I(seg_16_28_sp4_h_r_2_67731),
    .O(seg_16_28_local_g0_2_67635)
  );
  Span4Mux_h4 t3139 (
    .I(seg_16_28_sp4_v_b_8_63548),
    .O(seg_16_28_sp4_h_r_2_67731)
  );
  CascadeMux t314 (
    .I(net_53759),
    .O(net_53759_cascademuxed)
  );
  LocalMux t3140 (
    .I(seg_16_28_neigh_op_top_0_63884),
    .O(seg_16_28_local_g0_0_67633)
  );
  LocalMux t3141 (
    .I(seg_16_29_lutff_2_out_63886),
    .O(seg_16_29_local_g2_2_67774)
  );
  LocalMux t3142 (
    .I(seg_16_28_neigh_op_top_4_63888),
    .O(seg_16_28_local_g0_4_67637)
  );
  LocalMux t3143 (
    .I(seg_16_29_lutff_6_out_63890),
    .O(seg_16_29_local_g2_6_67778)
  );
  LocalMux t3144 (
    .I(seg_17_9_sp12_v_b_0_68077),
    .O(seg_17_9_local_g3_0_69151)
  );
  LocalMux t3145 (
    .I(seg_16_9_sp4_r_v_b_17_65161),
    .O(seg_16_9_local_g3_1_65321)
  );
  Span4Mux_v4 t3146 (
    .I(seg_17_6_sp4_v_b_8_64673),
    .O(seg_16_9_sp4_r_v_b_17_65161)
  );
  Span4Mux_v4 t3147 (
    .I(seg_17_2_sp4_v_b_5_64390),
    .O(seg_17_6_sp4_v_b_8_64673)
  );
  LocalMux t3148 (
    .I(seg_16_9_sp4_r_v_b_14_65158),
    .O(seg_16_9_local_g2_6_65318)
  );
  Span4Mux_v4 t3149 (
    .I(seg_17_6_sp4_v_b_3_64666),
    .O(seg_16_9_sp4_r_v_b_14_65158)
  );
  Span4Mux_v4 t3150 (
    .I(seg_17_2_sp4_v_b_7_64392),
    .O(seg_17_6_sp4_v_b_3_64666)
  );
  LocalMux t3151 (
    .I(seg_16_5_neigh_op_rgt_0_64763),
    .O(seg_16_5_local_g2_0_64820)
  );
  LocalMux t3152 (
    .I(seg_17_5_lutff_0_out_64763),
    .O(seg_17_5_local_g3_0_68659)
  );
  LocalMux t3153 (
    .I(seg_16_5_neigh_op_rgt_1_64764),
    .O(seg_16_5_local_g3_1_64829)
  );
  LocalMux t3154 (
    .I(seg_17_6_neigh_op_bot_1_64764),
    .O(seg_17_6_local_g0_1_68759)
  );
  LocalMux t3155 (
    .I(seg_16_5_neigh_op_rgt_2_64765),
    .O(seg_16_5_local_g3_2_64830)
  );
  LocalMux t3156 (
    .I(seg_17_6_neigh_op_bot_2_64765),
    .O(seg_17_6_local_g1_2_68768)
  );
  LocalMux t3157 (
    .I(seg_16_5_neigh_op_rgt_3_64766),
    .O(seg_16_5_local_g3_3_64831)
  );
  LocalMux t3158 (
    .I(seg_17_5_lutff_3_out_64766),
    .O(seg_17_5_local_g3_3_68662)
  );
  LocalMux t3159 (
    .I(seg_18_6_neigh_op_bnl_5_64768),
    .O(seg_18_6_local_g2_5_72610)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t316 (
    .carryinitin(),
    .carryinitout(t315)
  );
  LocalMux t3160 (
    .I(seg_16_5_neigh_op_rgt_6_64769),
    .O(seg_16_5_local_g3_6_64834)
  );
  LocalMux t3161 (
    .I(seg_17_6_neigh_op_bot_6_64769),
    .O(seg_17_6_local_g0_6_68764)
  );
  LocalMux t3162 (
    .I(seg_16_5_neigh_op_rgt_7_64770),
    .O(seg_16_5_local_g2_7_64827)
  );
  LocalMux t3163 (
    .I(seg_17_5_lutff_7_out_64770),
    .O(seg_17_5_local_g3_7_68666)
  );
  LocalMux t3164 (
    .I(seg_17_6_neigh_op_bot_7_64770),
    .O(seg_17_6_local_g1_7_68773)
  );
  LocalMux t3165 (
    .I(seg_16_6_neigh_op_rgt_0_64886),
    .O(seg_16_6_local_g2_0_64943)
  );
  LocalMux t3166 (
    .I(seg_17_6_lutff_0_out_64886),
    .O(seg_17_6_local_g0_0_68758)
  );
  LocalMux t3167 (
    .I(seg_17_6_lutff_0_out_64886),
    .O(seg_17_6_local_g2_0_68774)
  );
  LocalMux t3168 (
    .I(seg_18_6_neigh_op_lft_4_64890),
    .O(seg_18_6_local_g1_4_72601)
  );
  LocalMux t3169 (
    .I(seg_18_6_neigh_op_lft_5_64891),
    .O(seg_18_6_local_g1_5_72602)
  );
  LocalMux t3170 (
    .I(seg_18_6_neigh_op_lft_7_64893),
    .O(seg_18_6_local_g1_7_72604)
  );
  LocalMux t3171 (
    .I(seg_16_10_neigh_op_bnr_1_65256),
    .O(seg_16_10_local_g1_1_65428)
  );
  LocalMux t3172 (
    .I(seg_17_14_sp4_v_b_23_65782),
    .O(seg_17_14_local_g0_7_69749)
  );
  Span4Mux_v4 t3173 (
    .I(seg_17_11_sp4_v_b_10_65290),
    .O(seg_17_14_sp4_v_b_23_65782)
  );
  LocalMux t3174 (
    .I(seg_20_13_sp4_v_b_42_77119),
    .O(seg_20_13_local_g2_2_80499)
  );
  Span4Mux_v4 t3175 (
    .I(seg_20_12_sp4_h_l_42_65768),
    .O(seg_20_13_sp4_v_b_42_77119)
  );
  LocalMux t3176 (
    .I(seg_18_13_neigh_op_lft_3_65750),
    .O(seg_18_13_local_g0_3_73453)
  );
  LocalMux t3177 (
    .I(seg_17_15_sp4_r_v_b_5_69606),
    .O(seg_17_15_local_g1_5_69878)
  );
  LocalMux t3178 (
    .I(seg_17_15_neigh_op_bot_0_65870),
    .O(seg_17_15_local_g1_0_69873)
  );
  LocalMux t3179 (
    .I(seg_18_14_neigh_op_lft_2_65872),
    .O(seg_18_14_local_g1_2_73583)
  );
  CascadeMux t318 (
    .I(net_53840),
    .O(net_53840_cascademuxed)
  );
  LocalMux t3180 (
    .I(seg_18_14_neigh_op_lft_3_65873),
    .O(seg_18_14_local_g0_3_73576)
  );
  LocalMux t3181 (
    .I(seg_18_14_neigh_op_lft_4_65874),
    .O(seg_18_14_local_g1_4_73585)
  );
  LocalMux t3182 (
    .I(seg_17_14_lutff_5_out_65875),
    .O(seg_17_14_local_g2_5_69763)
  );
  LocalMux t3183 (
    .I(seg_18_14_neigh_op_lft_7_65877),
    .O(seg_18_14_local_g0_7_73580)
  );
  LocalMux t3184 (
    .I(seg_19_16_sp4_h_r_14_73918),
    .O(seg_19_16_local_g0_6_77339)
  );
  Span4Mux_h4 t3185 (
    .I(seg_18_16_sp4_v_b_3_69727),
    .O(seg_19_16_sp4_h_r_14_73918)
  );
  LocalMux t3186 (
    .I(seg_17_14_neigh_op_top_0_65993),
    .O(seg_17_14_local_g0_0_69742)
  );
  LocalMux t3187 (
    .I(seg_17_15_lutff_4_out_65997),
    .O(seg_17_15_local_g1_4_69877)
  );
  LocalMux t3188 (
    .I(seg_21_15_sp4_h_r_9_84663),
    .O(seg_21_15_local_g1_1_84567)
  );
  Span4Mux_h4 t3189 (
    .I(seg_21_15_sp4_h_l_43_69967),
    .O(seg_21_15_sp4_h_r_9_84663)
  );
  CascadeMux t319 (
    .I(net_53846),
    .O(net_53846_cascademuxed)
  );
  LocalMux t3190 (
    .I(seg_17_17_neigh_op_bot_1_66117),
    .O(seg_17_17_local_g0_1_70112)
  );
  LocalMux t3191 (
    .I(seg_13_16_sp4_h_r_22_50932),
    .O(seg_13_16_local_g0_6_54672)
  );
  Span4Mux_h4 t3192 (
    .I(seg_16_16_sp4_h_r_3_66256),
    .O(seg_13_16_sp4_h_r_22_50932)
  );
  LocalMux t3193 (
    .I(seg_15_16_sp4_h_r_6_62428),
    .O(seg_15_16_local_g1_6_62340)
  );
  LocalMux t3194 (
    .I(seg_18_17_neigh_op_lft_0_66239),
    .O(seg_18_17_local_g1_0_73950)
  );
  LocalMux t3195 (
    .I(seg_17_17_lutff_2_out_66241),
    .O(seg_17_17_local_g3_2_70137)
  );
  LocalMux t3196 (
    .I(seg_19_17_sp4_h_r_34_70207),
    .O(seg_19_17_local_g2_2_77453)
  );
  LocalMux t3197 (
    .I(seg_20_17_sp4_h_r_3_81072),
    .O(seg_20_17_local_g1_3_80984)
  );
  Span4Mux_h4 t3198 (
    .I(seg_20_17_sp4_h_l_38_66379),
    .O(seg_20_17_sp4_h_r_3_81072)
  );
  LocalMux t3199 (
    .I(seg_19_17_sp4_h_r_26_70209),
    .O(seg_19_17_local_g3_2_77461)
  );
  CascadeMux t32 (
    .I(net_17526),
    .O(net_17526_cascademuxed)
  );
  CascadeMux t320 (
    .I(net_53852),
    .O(net_53852_cascademuxed)
  );
  LocalMux t3200 (
    .I(seg_18_18_neigh_op_lft_0_66362),
    .O(seg_18_18_local_g0_0_74065)
  );
  LocalMux t3201 (
    .I(seg_18_18_neigh_op_lft_1_66363),
    .O(seg_18_18_local_g1_1_74074)
  );
  LocalMux t3202 (
    .I(seg_17_17_neigh_op_top_2_66364),
    .O(seg_17_17_local_g0_2_70113)
  );
  LocalMux t3203 (
    .I(seg_18_18_neigh_op_lft_4_66366),
    .O(seg_18_18_local_g1_4_74077)
  );
  LocalMux t3204 (
    .I(seg_15_27_sp12_v_b_7_62665),
    .O(seg_15_27_local_g3_7_63710)
  );
  Span12Mux_v12 t3205 (
    .I(seg_15_18_sp12_h_r_0_62662),
    .O(seg_15_27_sp12_v_b_7_62665)
  );
  LocalMux t3206 (
    .I(seg_15_28_sp12_v_b_4_62665),
    .O(seg_15_28_local_g3_4_63830)
  );
  Span12Mux_v12 t3207 (
    .I(seg_15_18_sp12_h_r_0_62662),
    .O(seg_15_28_sp12_v_b_4_62665)
  );
  LocalMux t3208 (
    .I(seg_16_29_sp4_v_b_18_63791),
    .O(seg_16_29_local_g0_2_67758)
  );
  Span4Mux_v4 t3209 (
    .I(seg_16_26_sp4_v_b_4_63298),
    .O(seg_16_29_sp4_v_b_18_63791)
  );
  CascadeMux t321 (
    .I(net_53870),
    .O(net_53870_cascademuxed)
  );
  Span4Mux_v4 t3210 (
    .I(seg_16_22_sp4_v_b_1_62801),
    .O(seg_16_26_sp4_v_b_4_63298)
  );
  Span4Mux_v4 t3211 (
    .I(seg_16_18_sp4_h_r_1_66498),
    .O(seg_16_22_sp4_v_b_1_62801)
  );
  LocalMux t3212 (
    .I(seg_18_18_sp4_h_r_27_66502),
    .O(seg_18_18_local_g2_3_74084)
  );
  LocalMux t3213 (
    .I(seg_20_18_sp4_h_r_11_81193),
    .O(seg_20_18_local_g1_3_81107)
  );
  Span4Mux_h4 t3214 (
    .I(seg_20_18_sp4_h_l_46_66500),
    .O(seg_20_18_sp4_h_r_11_81193)
  );
  LocalMux t3215 (
    .I(seg_14_26_sp4_v_b_11_55643),
    .O(seg_14_26_local_g1_3_59737)
  );
  Span4Mux_v4 t3216 (
    .I(seg_14_22_sp4_v_b_3_55143),
    .O(seg_14_26_sp4_v_b_11_55643)
  );
  Span4Mux_v4 t3217 (
    .I(seg_14_18_sp4_h_r_9_58847),
    .O(seg_14_22_sp4_v_b_3_55143)
  );
  LocalMux t3218 (
    .I(seg_14_28_sp4_v_b_20_56010),
    .O(seg_14_28_local_g1_4_59984)
  );
  Span4Mux_v4 t3219 (
    .I(seg_14_25_sp4_h_r_9_59708),
    .O(seg_14_28_sp4_v_b_20_56010)
  );
  CascadeMux t322 (
    .I(net_53876),
    .O(net_53876_cascademuxed)
  );
  Span4Mux_h4 t3220 (
    .I(seg_18_25_sp4_v_b_4_70837),
    .O(seg_14_25_sp4_h_r_9_59708)
  );
  Span4Mux_v4 t3221 (
    .I(seg_18_21_sp4_v_b_8_70349),
    .O(seg_18_25_sp4_v_b_4_70837)
  );
  LocalMux t3222 (
    .I(seg_16_28_sp4_r_v_b_16_67497),
    .O(seg_16_28_local_g3_0_67657)
  );
  Span4Mux_v4 t3223 (
    .I(seg_17_25_sp4_v_b_9_67009),
    .O(seg_16_28_sp4_r_v_b_16_67497)
  );
  Span4Mux_v4 t3224 (
    .I(seg_17_21_sp4_v_b_9_66517),
    .O(seg_17_25_sp4_v_b_9_67009)
  );
  LocalMux t3225 (
    .I(seg_17_19_lutff_1_out_66486),
    .O(seg_17_19_local_g2_1_70374)
  );
  LocalMux t3226 (
    .I(seg_17_19_lutff_5_out_66490),
    .O(seg_17_19_local_g0_5_70362)
  );
  LocalMux t3227 (
    .I(seg_17_18_neigh_op_top_6_66491),
    .O(seg_17_18_local_g1_6_70248)
  );
  LocalMux t3228 (
    .I(seg_17_19_lutff_7_out_66492),
    .O(seg_17_19_local_g3_7_70388)
  );
  LocalMux t3229 (
    .I(seg_19_18_sp4_v_b_19_73932),
    .O(seg_19_18_local_g1_3_77548)
  );
  CascadeMux t323 (
    .I(net_54209),
    .O(net_54209_cascademuxed)
  );
  Span4Mux_v4 t3230 (
    .I(seg_19_19_sp4_h_l_37_62789),
    .O(seg_19_18_sp4_v_b_19_73932)
  );
  LocalMux t3231 (
    .I(seg_20_19_sp4_h_r_45_70461),
    .O(seg_20_19_local_g2_5_81240)
  );
  LocalMux t3232 (
    .I(seg_19_17_sp4_h_r_16_74043),
    .O(seg_19_17_local_g0_0_77435)
  );
  Span4Mux_h4 t3233 (
    .I(seg_18_17_sp4_v_t_40_70344),
    .O(seg_19_17_sp4_h_r_16_74043)
  );
  LocalMux t3234 (
    .I(seg_17_19_neigh_op_top_0_66608),
    .O(seg_17_19_local_g1_0_70365)
  );
  LocalMux t3235 (
    .I(seg_18_20_neigh_op_lft_1_66609),
    .O(seg_18_20_local_g1_1_74320)
  );
  LocalMux t3236 (
    .I(seg_16_20_neigh_op_rgt_2_66610),
    .O(seg_16_20_local_g3_2_66675)
  );
  LocalMux t3237 (
    .I(seg_17_20_lutff_5_out_66613),
    .O(seg_17_20_local_g2_5_70501)
  );
  LocalMux t3238 (
    .I(seg_17_20_lutff_6_out_66614),
    .O(seg_17_20_local_g2_6_70502)
  );
  LocalMux t3239 (
    .I(seg_19_17_sp4_h_r_31_70214),
    .O(seg_19_17_local_g3_7_77466)
  );
  CascadeMux t324 (
    .I(net_54215),
    .O(net_54215_cascademuxed)
  );
  Span4Mux_h4 t3240 (
    .I(seg_17_17_sp4_v_t_42_66515),
    .O(seg_19_17_sp4_h_r_31_70214)
  );
  LocalMux t3241 (
    .I(seg_17_20_neigh_op_top_6_66737),
    .O(seg_17_20_local_g1_6_70494)
  );
  LocalMux t3242 (
    .I(seg_17_15_sp4_r_v_b_31_69854),
    .O(seg_17_15_local_g1_7_69880)
  );
  Span4Mux_v4 t3243 (
    .I(seg_18_17_sp4_v_t_46_70350),
    .O(seg_17_15_sp4_r_v_b_31_69854)
  );
  LocalMux t3244 (
    .I(seg_17_16_sp4_r_v_b_18_69854),
    .O(seg_17_16_local_g3_2_70014)
  );
  Span4Mux_v4 t3245 (
    .I(seg_18_17_sp4_v_t_46_70350),
    .O(seg_17_16_sp4_r_v_b_18_69854)
  );
  LocalMux t3246 (
    .I(seg_18_31_span4_vert_5_71574),
    .O(seg_18_31_local_g0_5_75682)
  );
  LocalMux t3247 (
    .I(seg_16_29_sp4_r_v_b_32_67748),
    .O(seg_16_29_local_g0_3_67759)
  );
  LocalMux t3248 (
    .I(seg_16_29_sp4_r_v_b_32_67748),
    .O(seg_16_29_local_g2_0_67772)
  );
  LocalMux t3249 (
    .I(seg_16_2_sp4_r_v_b_12_64400),
    .O(seg_16_2_local_g2_4_64455)
  );
  CascadeMux t325 (
    .I(net_54221),
    .O(net_54221_cascademuxed)
  );
  IoSpan4Mux t3250 (
    .I(seg_17_0_span4_horz_r_0_68093),
    .O(seg_16_2_sp4_r_v_b_12_64400)
  );
  LocalMux t3251 (
    .I(seg_17_6_neigh_op_bnr_5_68599),
    .O(seg_17_6_local_g1_5_68771)
  );
  LocalMux t3252 (
    .I(seg_18_5_lutff_5_out_68599),
    .O(seg_18_5_local_g3_5_72495)
  );
  LocalMux t3253 (
    .I(seg_18_6_neigh_op_bot_5_68599),
    .O(seg_18_6_local_g0_5_72594)
  );
  LocalMux t3254 (
    .I(seg_18_5_lutff_7_out_68601),
    .O(seg_18_5_local_g3_7_72497)
  );
  LocalMux t3255 (
    .I(seg_16_5_sp4_h_r_18_61076),
    .O(seg_16_5_local_g1_2_64814)
  );
  LocalMux t3256 (
    .I(seg_17_5_neigh_op_tnr_0_68717),
    .O(seg_17_5_local_g2_0_68651)
  );
  LocalMux t3257 (
    .I(seg_17_6_neigh_op_rgt_0_68717),
    .O(seg_17_6_local_g3_0_68782)
  );
  LocalMux t3258 (
    .I(seg_18_5_neigh_op_top_0_68717),
    .O(seg_18_5_local_g0_0_72466)
  );
  LocalMux t3259 (
    .I(seg_18_6_lutff_0_out_68717),
    .O(seg_18_6_local_g1_0_72597)
  );
  CascadeMux t326 (
    .I(net_54227),
    .O(net_54227_cascademuxed)
  );
  LocalMux t3260 (
    .I(seg_18_6_lutff_2_out_68719),
    .O(seg_18_6_local_g2_2_72607)
  );
  LocalMux t3261 (
    .I(seg_18_6_lutff_5_out_68722),
    .O(seg_18_6_local_g3_5_72618)
  );
  LocalMux t3262 (
    .I(seg_17_6_neigh_op_rgt_7_68724),
    .O(seg_17_6_local_g2_7_68781)
  );
  LocalMux t3263 (
    .I(seg_18_6_lutff_7_out_68724),
    .O(seg_18_6_local_g2_7_72612)
  );
  LocalMux t3264 (
    .I(seg_20_6_sp4_h_r_34_72685),
    .O(seg_20_6_local_g2_2_79638)
  );
  LocalMux t3265 (
    .I(seg_20_6_sp4_h_r_26_72687),
    .O(seg_20_6_local_g3_2_79646)
  );
  LocalMux t3266 (
    .I(seg_21_9_sp4_r_v_b_15_83683),
    .O(seg_21_9_local_g2_7_83843)
  );
  Span4Mux_v4 t3267 (
    .I(seg_22_6_sp4_h_l_39_72687),
    .O(seg_21_9_sp4_r_v_b_15_83683)
  );
  LocalMux t3268 (
    .I(seg_16_5_sp4_v_b_22_60843),
    .O(seg_16_5_local_g1_6_64818)
  );
  Span4Mux_v4 t3269 (
    .I(seg_16_6_sp4_h_r_6_65029),
    .O(seg_16_5_sp4_v_b_22_60843)
  );
  CascadeMux t327 (
    .I(net_54245),
    .O(net_54245_cascademuxed)
  );
  LocalMux t3270 (
    .I(seg_18_6_sp4_r_v_b_3_72328),
    .O(seg_18_6_local_g1_3_72600)
  );
  Span4Mux_v4 t3271 (
    .I(seg_19_6_sp4_h_l_44_61201),
    .O(seg_18_6_sp4_r_v_b_3_72328)
  );
  LocalMux t3272 (
    .I(seg_12_8_sp4_r_v_b_31_49840),
    .O(seg_12_8_local_g1_7_49866)
  );
  Span4Mux_v4 t3273 (
    .I(seg_13_10_sp4_h_r_2_54026),
    .O(seg_12_8_sp4_r_v_b_31_49840)
  );
  Span4Mux_h4 t3274 (
    .I(seg_17_10_sp4_h_r_11_69347),
    .O(seg_13_10_sp4_h_r_2_54026)
  );
  LocalMux t3275 (
    .I(seg_13_9_sp4_v_b_18_49840),
    .O(seg_13_9_local_g1_2_53815)
  );
  Span4Mux_v4 t3276 (
    .I(seg_13_10_sp4_h_r_2_54026),
    .O(seg_13_9_sp4_v_b_18_49840)
  );
  LocalMux t3277 (
    .I(seg_10_8_sp4_r_v_b_32_42181),
    .O(seg_10_8_local_g0_3_42192)
  );
  Span4Mux_v4 t3278 (
    .I(seg_11_10_sp4_h_r_3_46365),
    .O(seg_10_8_sp4_r_v_b_32_42181)
  );
  Span4Mux_h4 t3279 (
    .I(seg_15_10_sp4_h_r_3_61687),
    .O(seg_11_10_sp4_h_r_3_46365)
  );
  CascadeMux t328 (
    .I(net_54332),
    .O(net_54332_cascademuxed)
  );
  LocalMux t3280 (
    .I(seg_10_8_sp4_r_v_b_30_42179),
    .O(seg_10_8_local_g0_6_42195)
  );
  Span4Mux_v4 t3281 (
    .I(seg_11_10_sp4_h_r_6_46368),
    .O(seg_10_8_sp4_r_v_b_30_42179)
  );
  Span4Mux_h4 t3282 (
    .I(seg_15_10_sp4_h_r_3_61687),
    .O(seg_11_10_sp4_h_r_6_46368)
  );
  LocalMux t3283 (
    .I(seg_11_7_sp4_v_b_43_42179),
    .O(seg_11_7_local_g3_3_45924)
  );
  Span4Mux_v4 t3284 (
    .I(seg_11_10_sp4_h_r_6_46368),
    .O(seg_11_7_sp4_v_b_43_42179)
  );
  LocalMux t3285 (
    .I(seg_11_9_sp4_v_b_14_42174),
    .O(seg_11_9_local_g1_6_46157)
  );
  Span4Mux_v4 t3286 (
    .I(seg_11_10_sp4_h_r_3_46365),
    .O(seg_11_9_sp4_v_b_14_42174)
  );
  LocalMux t3287 (
    .I(seg_14_7_sp4_r_v_b_45_57504),
    .O(seg_14_7_local_g3_5_57418)
  );
  Span4Mux_v4 t3288 (
    .I(seg_15_10_sp4_h_r_3_61687),
    .O(seg_14_7_sp4_r_v_b_45_57504)
  );
  LocalMux t3289 (
    .I(seg_14_8_sp4_r_v_b_32_57504),
    .O(seg_14_8_local_g2_0_57528)
  );
  CascadeMux t329 (
    .I(net_54338),
    .O(net_54338_cascademuxed)
  );
  Span4Mux_v4 t3290 (
    .I(seg_15_10_sp4_h_r_3_61687),
    .O(seg_14_8_sp4_r_v_b_32_57504)
  );
  LocalMux t3291 (
    .I(seg_21_16_sp4_r_v_b_33_84672),
    .O(seg_21_16_local_g2_1_84698)
  );
  Span4Mux_v4 t3292 (
    .I(seg_22_14_sp4_v_b_6_84179),
    .O(seg_21_16_sp4_r_v_b_33_84672)
  );
  Span4Mux_v4 t3293 (
    .I(seg_22_10_sp4_h_l_43_73183),
    .O(seg_22_14_sp4_v_b_6_84179)
  );
  LocalMux t3294 (
    .I(seg_22_17_sp4_v_b_15_84667),
    .O(seg_22_17_local_g1_7_88650)
  );
  Span4Mux_v4 t3295 (
    .I(seg_22_14_sp4_v_b_6_84179),
    .O(seg_22_17_sp4_v_b_15_84667)
  );
  LocalMux t3296 (
    .I(seg_10_7_sp4_h_r_5_42167),
    .O(seg_10_7_local_g0_5_42071)
  );
  Span4Mux_h4 t3297 (
    .I(seg_14_7_sp4_h_r_5_57490),
    .O(seg_10_7_sp4_h_r_5_42167)
  );
  Span4Mux_h4 t3298 (
    .I(seg_18_7_sp4_v_t_46_69120),
    .O(seg_14_7_sp4_h_r_5_57490)
  );
  LocalMux t3299 (
    .I(seg_20_12_sp4_h_r_36_69591),
    .O(seg_20_12_local_g2_4_80378)
  );
  CascadeMux t33 (
    .I(net_17544),
    .O(net_17544_cascademuxed)
  );
  CascadeMux t330 (
    .I(net_54344),
    .O(net_54344_cascademuxed)
  );
  LocalMux t3300 (
    .I(seg_20_12_sp4_h_r_2_80456),
    .O(seg_20_12_local_g0_2_80360)
  );
  Span4Mux_h4 t3301 (
    .I(seg_20_12_sp4_h_l_43_65767),
    .O(seg_20_12_sp4_h_r_2_80456)
  );
  LocalMux t3302 (
    .I(seg_20_12_sp4_h_r_30_73429),
    .O(seg_20_12_local_g2_6_80380)
  );
  LocalMux t3303 (
    .I(seg_18_14_neigh_op_bot_1_69579),
    .O(seg_18_14_local_g1_1_73582)
  );
  LocalMux t3304 (
    .I(seg_20_13_sp12_h_r_8_65878),
    .O(seg_20_13_local_g0_0_80481)
  );
  LocalMux t3305 (
    .I(seg_21_13_sp4_h_r_37_73544),
    .O(seg_21_13_local_g3_5_84341)
  );
  LocalMux t3306 (
    .I(seg_20_13_sp4_h_r_38_69718),
    .O(seg_20_13_local_g2_6_80503)
  );
  LocalMux t3307 (
    .I(seg_21_15_sp4_v_b_28_80715),
    .O(seg_21_15_local_g3_4_84586)
  );
  Span4Mux_v4 t3308 (
    .I(seg_21_13_sp4_h_l_46_69716),
    .O(seg_21_15_sp4_v_b_28_80715)
  );
  LocalMux t3309 (
    .I(seg_21_13_sp4_h_r_23_80577),
    .O(seg_21_13_local_g1_7_84327)
  );
  CascadeMux t331 (
    .I(net_54356),
    .O(net_54356_cascademuxed)
  );
  Span4Mux_h4 t3310 (
    .I(seg_20_13_sp4_h_l_39_65886),
    .O(seg_21_13_sp4_h_r_23_80577)
  );
  LocalMux t3311 (
    .I(seg_20_13_sp4_h_r_28_73550),
    .O(seg_20_13_local_g3_4_80509)
  );
  LocalMux t3312 (
    .I(seg_21_13_sp4_h_r_45_73554),
    .O(seg_21_13_local_g2_5_84333)
  );
  LocalMux t3313 (
    .I(seg_18_14_lutff_1_out_69702),
    .O(seg_18_14_local_g2_1_73590)
  );
  LocalMux t3314 (
    .I(seg_18_13_neigh_op_top_4_69705),
    .O(seg_18_13_local_g0_4_73454)
  );
  LocalMux t3315 (
    .I(seg_18_14_lutff_7_out_69708),
    .O(seg_18_14_local_g2_7_73596)
  );
  LocalMux t3316 (
    .I(seg_20_14_sp4_h_r_24_73667),
    .O(seg_20_14_local_g2_0_80620)
  );
  LocalMux t3317 (
    .I(seg_20_14_sp4_h_r_34_73669),
    .O(seg_20_14_local_g2_2_80622)
  );
  LocalMux t3318 (
    .I(seg_20_14_sp4_h_r_44_69847),
    .O(seg_20_14_local_g2_4_80624)
  );
  LocalMux t3319 (
    .I(seg_20_14_sp4_h_r_30_73675),
    .O(seg_20_14_local_g2_6_80626)
  );
  CascadeMux t332 (
    .I(net_54374),
    .O(net_54374_cascademuxed)
  );
  LocalMux t3320 (
    .I(seg_20_15_sp4_h_r_24_73790),
    .O(seg_20_15_local_g3_0_80751)
  );
  LocalMux t3321 (
    .I(seg_20_15_sp4_h_r_38_69964),
    .O(seg_20_15_local_g2_6_80749)
  );
  LocalMux t3322 (
    .I(seg_20_15_sp4_h_r_44_69970),
    .O(seg_20_15_local_g2_4_80747)
  );
  LocalMux t3323 (
    .I(seg_20_15_sp4_h_r_21_77315),
    .O(seg_20_15_local_g1_5_80740)
  );
  Span4Mux_h4 t3324 (
    .I(seg_19_15_sp4_h_l_40_62304),
    .O(seg_20_15_sp4_h_r_21_77315)
  );
  LocalMux t3325 (
    .I(seg_20_15_sp4_h_r_16_77312),
    .O(seg_20_15_local_g1_0_80735)
  );
  Span4Mux_h4 t3326 (
    .I(seg_19_15_sp4_h_l_44_62308),
    .O(seg_20_15_sp4_h_r_16_77312)
  );
  LocalMux t3327 (
    .I(seg_20_15_sp4_h_r_22_77308),
    .O(seg_20_15_local_g1_6_80741)
  );
  Span4Mux_h4 t3328 (
    .I(seg_19_15_sp4_v_b_11_73443),
    .O(seg_20_15_sp4_h_r_22_77308)
  );
  LocalMux t3329 (
    .I(seg_20_15_sp4_h_r_18_77314),
    .O(seg_20_15_local_g0_2_80729)
  );
  CascadeMux t333 (
    .I(net_54455),
    .O(net_54455_cascademuxed)
  );
  Span4Mux_h4 t3330 (
    .I(seg_19_15_sp4_v_b_7_73439),
    .O(seg_20_15_sp4_h_r_18_77314)
  );
  LocalMux t3331 (
    .I(seg_18_16_lutff_2_out_69949),
    .O(seg_18_16_local_g3_2_73845)
  );
  LocalMux t3332 (
    .I(seg_19_16_neigh_op_lft_2_69949),
    .O(seg_19_16_local_g1_2_77343)
  );
  LocalMux t3333 (
    .I(seg_21_17_sp4_v_b_44_81087),
    .O(seg_21_17_local_g3_4_84832)
  );
  Span4Mux_v4 t3334 (
    .I(seg_21_16_sp4_h_l_44_70093),
    .O(seg_21_17_sp4_v_b_44_81087)
  );
  LocalMux t3335 (
    .I(seg_20_16_sp4_h_r_28_73919),
    .O(seg_20_16_local_g2_4_80870)
  );
  LocalMux t3336 (
    .I(seg_19_18_sp4_v_b_13_73926),
    .O(seg_19_18_local_g0_5_77542)
  );
  LocalMux t3337 (
    .I(seg_19_14_sp4_v_b_29_73560),
    .O(seg_19_14_local_g2_5_77150)
  );
  LocalMux t3338 (
    .I(seg_21_17_sp4_h_r_37_74036),
    .O(seg_21_17_local_g2_5_84825)
  );
  LocalMux t3339 (
    .I(seg_22_17_sp4_h_r_3_88734),
    .O(seg_22_17_local_g1_3_88646)
  );
  CascadeMux t334 (
    .I(net_54461),
    .O(net_54461_cascademuxed)
  );
  Span4Mux_h4 t3340 (
    .I(seg_22_17_sp4_h_l_37_74036),
    .O(seg_22_17_sp4_h_r_3_88734)
  );
  LocalMux t3341 (
    .I(seg_21_14_sp4_r_v_b_47_84552),
    .O(seg_21_14_local_g3_7_84466)
  );
  Span4Mux_v4 t3342 (
    .I(seg_22_17_sp4_h_l_47_74038),
    .O(seg_21_14_sp4_r_v_b_47_84552)
  );
  LocalMux t3343 (
    .I(seg_20_17_sp4_h_r_36_70206),
    .O(seg_20_17_local_g2_4_80993)
  );
  LocalMux t3344 (
    .I(seg_22_17_sp4_h_r_17_84904),
    .O(seg_22_17_local_g0_1_88636)
  );
  Span4Mux_h4 t3345 (
    .I(seg_21_17_sp4_h_l_36_70206),
    .O(seg_22_17_sp4_h_r_17_84904)
  );
  LocalMux t3346 (
    .I(seg_20_17_sp4_h_r_26_74040),
    .O(seg_20_17_local_g2_2_80991)
  );
  LocalMux t3347 (
    .I(seg_20_17_sp4_h_r_2_81071),
    .O(seg_20_17_local_g0_2_80975)
  );
  Span4Mux_h4 t3348 (
    .I(seg_20_17_sp4_h_l_43_66382),
    .O(seg_20_17_sp4_h_r_2_81071)
  );
  LocalMux t3349 (
    .I(seg_20_17_sp4_h_r_19_77517),
    .O(seg_20_17_local_g0_3_80976)
  );
  CascadeMux t335 (
    .I(net_54467),
    .O(net_54467_cascademuxed)
  );
  Span4Mux_h4 t3350 (
    .I(seg_19_17_sp4_h_l_38_62548),
    .O(seg_20_17_sp4_h_r_19_77517)
  );
  LocalMux t3351 (
    .I(seg_21_17_sp4_h_r_41_74042),
    .O(seg_21_17_local_g2_1_84821)
  );
  LocalMux t3352 (
    .I(seg_22_17_sp4_h_r_4_88735),
    .O(seg_22_17_local_g1_4_88647)
  );
  Span4Mux_h4 t3353 (
    .I(seg_22_17_sp4_h_l_41_74042),
    .O(seg_22_17_sp4_h_r_4_88735)
  );
  LocalMux t3354 (
    .I(seg_20_17_sp4_h_r_32_74046),
    .O(seg_20_17_local_g3_0_80997)
  );
  LocalMux t3355 (
    .I(seg_18_18_lutff_3_out_70196),
    .O(seg_18_18_local_g3_3_74092)
  );
  LocalMux t3356 (
    .I(seg_18_17_neigh_op_top_4_70197),
    .O(seg_18_17_local_g0_4_73946)
  );
  LocalMux t3357 (
    .I(seg_18_18_lutff_5_out_70198),
    .O(seg_18_18_local_g0_5_74070)
  );
  LocalMux t3358 (
    .I(seg_21_18_sp4_h_r_4_85027),
    .O(seg_21_18_local_g0_4_84931)
  );
  Span4Mux_h4 t3359 (
    .I(seg_21_18_sp4_h_l_36_70329),
    .O(seg_21_18_sp4_h_r_4_85027)
  );
  CascadeMux t336 (
    .I(net_54473),
    .O(net_54473_cascademuxed)
  );
  LocalMux t3360 (
    .I(seg_20_18_sp4_h_r_9_81201),
    .O(seg_20_18_local_g1_1_81105)
  );
  Span4Mux_h4 t3361 (
    .I(seg_20_18_sp4_h_l_43_66505),
    .O(seg_20_18_sp4_h_r_9_81201)
  );
  LocalMux t3362 (
    .I(seg_21_18_sp4_h_r_41_74165),
    .O(seg_21_18_local_g3_1_84952)
  );
  LocalMux t3363 (
    .I(seg_18_18_neigh_op_top_7_70323),
    .O(seg_18_18_local_g1_7_74080)
  );
  LocalMux t3364 (
    .I(seg_20_18_sp4_h_r_18_77620),
    .O(seg_20_18_local_g0_2_81098)
  );
  Span4Mux_h4 t3365 (
    .I(seg_19_18_sp4_v_t_42_74300),
    .O(seg_20_18_sp4_h_r_18_77620)
  );
  LocalMux t3366 (
    .I(seg_15_22_sp4_h_r_23_59330),
    .O(seg_15_22_local_g1_7_63079)
  );
  Span4Mux_h4 t3367 (
    .I(seg_18_22_sp4_v_t_41_70960),
    .O(seg_15_22_sp4_h_r_23_59330)
  );
  Span4Mux_v4 t3368 (
    .I(seg_18_26_sp4_v_t_36_71447),
    .O(seg_18_22_sp4_v_t_41_70960)
  );
  Span4Mux_v4 t3369 (
    .I(seg_18_30_sp4_v_t_36_75655),
    .O(seg_18_26_sp4_v_t_36_71447)
  );
  CascadeMux t337 (
    .I(net_54491),
    .O(net_54491_cascademuxed)
  );
  LocalMux t3370 (
    .I(seg_15_23_sp4_h_r_12_59452),
    .O(seg_15_23_local_g0_4_63191)
  );
  Span4Mux_h4 t3371 (
    .I(seg_18_23_sp4_v_t_42_71084),
    .O(seg_15_23_sp4_h_r_12_59452)
  );
  Span4Mux_v4 t3372 (
    .I(seg_18_27_sp4_v_t_41_71575),
    .O(seg_18_23_sp4_v_t_42_71084)
  );
  LocalMux t3373 (
    .I(seg_17_21_sp4_r_v_b_27_70588),
    .O(seg_17_21_local_g0_3_70606)
  );
  Span4Mux_v4 t3374 (
    .I(seg_18_23_sp4_v_t_42_71084),
    .O(seg_17_21_sp4_r_v_b_27_70588)
  );
  LocalMux t3375 (
    .I(seg_15_23_sp4_h_r_13_59451),
    .O(seg_15_23_local_g0_5_63192)
  );
  Span4Mux_h4 t3376 (
    .I(seg_18_23_sp4_v_t_43_71085),
    .O(seg_15_23_sp4_h_r_13_59451)
  );
  Span4Mux_v4 t3377 (
    .I(seg_18_27_sp4_v_t_43_71577),
    .O(seg_18_23_sp4_v_t_43_71085)
  );
  LocalMux t3378 (
    .I(seg_20_13_neigh_op_lft_5_73414),
    .O(seg_20_13_local_g0_5_80486)
  );
  LocalMux t3379 (
    .I(seg_20_12_neigh_op_tnl_3_73412),
    .O(seg_20_12_local_g2_3_80377)
  );
  CascadeMux t338 (
    .I(net_54578),
    .O(net_54578_cascademuxed)
  );
  LocalMux t3380 (
    .I(seg_20_13_neigh_op_lft_2_73411),
    .O(seg_20_13_local_g1_2_80491)
  );
  LocalMux t3381 (
    .I(seg_18_14_neigh_op_bnr_1_73410),
    .O(seg_18_14_local_g0_1_73574)
  );
  LocalMux t3382 (
    .I(seg_18_14_neigh_op_bnr_7_73416),
    .O(seg_18_14_local_g1_7_73588)
  );
  LocalMux t3383 (
    .I(seg_21_13_sp4_h_r_24_77101),
    .O(seg_21_13_local_g2_0_84328)
  );
  LocalMux t3384 (
    .I(seg_17_13_sp4_h_r_0_69713),
    .O(seg_17_13_local_g1_0_69627)
  );
  LocalMux t3385 (
    .I(seg_17_13_sp4_h_r_20_65893),
    .O(seg_17_13_local_g0_4_69623)
  );
  LocalMux t3386 (
    .I(seg_20_13_neigh_op_tnl_6_73538),
    .O(seg_20_13_local_g3_6_80511)
  );
  LocalMux t3387 (
    .I(seg_20_13_neigh_op_tnl_5_73537),
    .O(seg_20_13_local_g3_5_80510)
  );
  LocalMux t3388 (
    .I(seg_20_13_neigh_op_tnl_2_73534),
    .O(seg_20_13_local_g3_2_80507)
  );
  LocalMux t3389 (
    .I(seg_21_13_sp4_r_v_b_22_84182),
    .O(seg_21_13_local_g3_6_84342)
  );
  CascadeMux t339 (
    .I(net_54596),
    .O(net_54596_cascademuxed)
  );
  Span4Mux_v4 t3390 (
    .I(seg_22_14_sp4_h_l_40_73674),
    .O(seg_21_13_sp4_r_v_b_22_84182)
  );
  LocalMux t3391 (
    .I(seg_20_12_sp4_v_b_27_76911),
    .O(seg_20_12_local_g3_3_80385)
  );
  LocalMux t3392 (
    .I(seg_21_13_sp4_h_r_17_80581),
    .O(seg_21_13_local_g0_1_84313)
  );
  Span4Mux_h4 t3393 (
    .I(seg_20_13_sp4_v_t_41_77220),
    .O(seg_21_13_sp4_h_r_17_80581)
  );
  LocalMux t3394 (
    .I(seg_21_13_sp4_h_r_14_80580),
    .O(seg_21_13_local_g1_6_84326)
  );
  Span4Mux_h4 t3395 (
    .I(seg_20_13_sp4_v_t_47_77226),
    .O(seg_21_13_sp4_h_r_14_80580)
  );
  LocalMux t3396 (
    .I(seg_20_12_sp4_v_b_31_76915),
    .O(seg_20_12_local_g2_7_80381)
  );
  LocalMux t3397 (
    .I(seg_18_14_neigh_op_tnr_5_73660),
    .O(seg_18_14_local_g3_5_73602)
  );
  LocalMux t3398 (
    .I(seg_20_15_neigh_op_lft_3_73658),
    .O(seg_20_15_local_g1_3_80738)
  );
  LocalMux t3399 (
    .I(seg_18_14_neigh_op_tnr_2_73657),
    .O(seg_18_14_local_g3_2_73599)
  );
  CascadeMux t34 (
    .I(net_20514),
    .O(net_20514_cascademuxed)
  );
  CascadeMux t340 (
    .I(net_54614),
    .O(net_54614_cascademuxed)
  );
  LocalMux t3400 (
    .I(seg_20_15_neigh_op_lft_1_73656),
    .O(seg_20_15_local_g1_1_80736)
  );
  LocalMux t3401 (
    .I(seg_20_15_neigh_op_lft_0_73655),
    .O(seg_20_15_local_g0_0_80727)
  );
  LocalMux t3402 (
    .I(seg_22_14_sp4_v_b_20_84303),
    .O(seg_22_14_local_g1_4_88278)
  );
  Span4Mux_v4 t3403 (
    .I(seg_22_15_sp4_h_l_38_73795),
    .O(seg_22_14_sp4_v_b_20_84303)
  );
  LocalMux t3404 (
    .I(seg_17_15_sp4_h_r_16_66135),
    .O(seg_17_15_local_g0_0_69865)
  );
  LocalMux t3405 (
    .I(seg_20_13_sp4_v_b_37_77114),
    .O(seg_20_13_local_g2_5_80502)
  );
  LocalMux t3406 (
    .I(seg_20_15_neigh_op_tnl_6_73784),
    .O(seg_20_15_local_g3_6_80757)
  );
  LocalMux t3407 (
    .I(seg_20_15_neigh_op_tnl_4_73782),
    .O(seg_20_15_local_g3_4_80755)
  );
  LocalMux t3408 (
    .I(seg_20_15_neigh_op_tnl_2_73780),
    .O(seg_20_15_local_g3_2_80753)
  );
  LocalMux t3409 (
    .I(seg_20_15_neigh_op_tnl_0_73778),
    .O(seg_20_15_local_g2_0_80743)
  );
  CascadeMux t341 (
    .I(net_54620),
    .O(net_54620_cascademuxed)
  );
  LocalMux t3410 (
    .I(seg_21_13_sp4_v_b_39_80590),
    .O(seg_21_13_local_g2_7_84335)
  );
  Span4Mux_v4 t3411 (
    .I(seg_21_16_sp4_h_l_39_70086),
    .O(seg_21_13_sp4_v_b_39_80590)
  );
  LocalMux t3412 (
    .I(seg_20_12_sp4_v_b_15_76810),
    .O(seg_20_12_local_g1_7_80373)
  );
  Span4Mux_v4 t3413 (
    .I(seg_20_13_sp4_v_t_43_77222),
    .O(seg_20_12_sp4_v_b_15_76810)
  );
  LocalMux t3414 (
    .I(seg_18_14_sp4_r_v_b_38_73681),
    .O(seg_18_14_local_g2_6_73595)
  );
  LocalMux t3415 (
    .I(seg_20_12_sp4_h_r_22_77002),
    .O(seg_20_12_local_g0_6_80364)
  );
  Span4Mux_h4 t3416 (
    .I(seg_19_12_sp4_v_t_43_73563),
    .O(seg_20_12_sp4_h_r_22_77002)
  );
  LocalMux t3417 (
    .I(seg_20_18_neigh_op_bnl_5_73906),
    .O(seg_20_18_local_g3_5_81125)
  );
  LocalMux t3418 (
    .I(seg_20_17_neigh_op_lft_4_73905),
    .O(seg_20_17_local_g1_4_80985)
  );
  LocalMux t3419 (
    .I(seg_20_18_neigh_op_bnl_3_73904),
    .O(seg_20_18_local_g2_3_81115)
  );
  CascadeMux t342 (
    .I(net_54701),
    .O(net_54701_cascademuxed)
  );
  LocalMux t3420 (
    .I(seg_18_18_neigh_op_bnr_7_73908),
    .O(seg_18_18_local_g0_7_74072)
  );
  LocalMux t3421 (
    .I(seg_22_16_sp4_r_v_b_19_88379),
    .O(seg_22_16_local_g3_3_88539)
  );
  Span4Mux_v4 t3422 (
    .I(seg_23_17_sp4_h_l_37_77509),
    .O(seg_22_16_sp4_r_v_b_19_88379)
  );
  LocalMux t3423 (
    .I(seg_17_17_sp4_h_r_29_62550),
    .O(seg_17_17_local_g3_5_70140)
  );
  Span4Mux_h4 t3424 (
    .I(seg_19_17_sp4_h_r_2_77513),
    .O(seg_17_17_sp4_h_r_29_62550)
  );
  LocalMux t3425 (
    .I(seg_20_17_sp4_h_r_41_70211),
    .O(seg_20_17_local_g3_1_80998)
  );
  LocalMux t3426 (
    .I(seg_20_13_sp4_v_b_8_76816),
    .O(seg_20_13_local_g1_0_80489)
  );
  Span4Mux_v4 t3427 (
    .I(seg_20_13_sp4_v_t_40_77219),
    .O(seg_20_13_sp4_v_b_8_76816)
  );
  LocalMux t3428 (
    .I(seg_20_18_neigh_op_lft_7_74031),
    .O(seg_20_18_local_g0_7_81103)
  );
  LocalMux t3429 (
    .I(seg_20_17_neigh_op_tnl_6_74030),
    .O(seg_20_17_local_g2_6_80995)
  );
  CascadeMux t343 (
    .I(net_54707),
    .O(net_54707_cascademuxed)
  );
  LocalMux t3430 (
    .I(seg_18_18_neigh_op_rgt_5_74029),
    .O(seg_18_18_local_g2_5_74086)
  );
  LocalMux t3431 (
    .I(seg_20_18_neigh_op_lft_3_74027),
    .O(seg_20_18_local_g0_3_81099)
  );
  LocalMux t3432 (
    .I(seg_18_18_neigh_op_rgt_2_74026),
    .O(seg_18_18_local_g3_2_74091)
  );
  LocalMux t3433 (
    .I(seg_18_18_neigh_op_rgt_1_74025),
    .O(seg_18_18_local_g2_1_74082)
  );
  LocalMux t3434 (
    .I(seg_20_17_neigh_op_tnl_0_74024),
    .O(seg_20_17_local_g2_0_80989)
  );
  LocalMux t3435 (
    .I(seg_17_17_sp4_h_r_35_62546),
    .O(seg_17_17_local_g3_3_70138)
  );
  Span4Mux_h4 t3436 (
    .I(seg_19_17_sp4_v_t_40_74175),
    .O(seg_17_17_sp4_h_r_35_62546)
  );
  LocalMux t3437 (
    .I(seg_20_6_lutff_2_out_76245),
    .O(seg_20_6_local_g1_2_79630)
  );
  LocalMux t3438 (
    .I(seg_20_6_lutff_5_out_76248),
    .O(seg_20_6_local_g2_5_79641)
  );
  LocalMux t3439 (
    .I(seg_21_6_neigh_op_lft_5_76248),
    .O(seg_21_6_local_g0_5_83456)
  );
  CascadeMux t344 (
    .I(net_54713),
    .O(net_54713_cascademuxed)
  );
  LocalMux t3440 (
    .I(seg_20_6_lutff_7_out_76250),
    .O(seg_20_6_local_g1_7_79635)
  );
  LocalMux t3441 (
    .I(seg_21_6_neigh_op_lft_7_76250),
    .O(seg_21_6_local_g1_7_83466)
  );
  LocalMux t3442 (
    .I(seg_18_6_sp4_h_r_24_65021),
    .O(seg_18_6_local_g2_0_72605)
  );
  Span4Mux_h4 t3443 (
    .I(seg_20_6_sp4_h_r_4_79720),
    .O(seg_18_6_sp4_h_r_24_65021)
  );
  LocalMux t3444 (
    .I(seg_20_6_sp4_r_v_b_33_79611),
    .O(seg_20_6_local_g0_2_79622)
  );
  LocalMux t3445 (
    .I(seg_20_6_neigh_op_top_0_76345),
    .O(seg_20_6_local_g1_0_79628)
  );
  LocalMux t3446 (
    .I(seg_18_6_sp4_r_v_b_16_72453),
    .O(seg_18_6_local_g3_0_72613)
  );
  Span4Mux_v4 t3447 (
    .I(seg_19_7_sp4_h_r_5_76496),
    .O(seg_18_6_sp4_r_v_b_16_72453)
  );
  LocalMux t3448 (
    .I(seg_17_6_sp4_v_b_19_64794),
    .O(seg_17_6_local_g1_3_68769)
  );
  Span4Mux_v4 t3449 (
    .I(seg_17_7_sp4_h_r_1_68976),
    .O(seg_17_6_sp4_v_b_19_64794)
  );
  CascadeMux t345 (
    .I(net_54719),
    .O(net_54719_cascademuxed)
  );
  Span4Mux_h4 t3450 (
    .I(seg_21_7_sp4_v_b_1_79480),
    .O(seg_17_7_sp4_h_r_1_68976)
  );
  LocalMux t3451 (
    .I(seg_17_5_sp4_h_r_3_68734),
    .O(seg_17_5_local_g1_3_68646)
  );
  Span4Mux_h4 t3452 (
    .I(seg_21_5_sp4_v_t_44_79734),
    .O(seg_17_5_sp4_h_r_3_68734)
  );
  LocalMux t3453 (
    .I(seg_18_5_sp4_h_r_26_64902),
    .O(seg_18_5_local_g2_2_72484)
  );
  Span4Mux_h4 t3454 (
    .I(seg_20_5_sp4_v_t_45_76408),
    .O(seg_18_5_sp4_h_r_26_64902)
  );
  LocalMux t3455 (
    .I(seg_20_9_lutff_1_out_76550),
    .O(seg_20_9_local_g3_1_80014)
  );
  LocalMux t3456 (
    .I(seg_20_10_neigh_op_bot_1_76550),
    .O(seg_20_10_local_g1_1_80121)
  );
  LocalMux t3457 (
    .I(seg_20_10_neigh_op_bot_5_76554),
    .O(seg_20_10_local_g0_5_80117)
  );
  LocalMux t3458 (
    .I(seg_21_9_neigh_op_lft_5_76554),
    .O(seg_21_9_local_g1_5_83833)
  );
  LocalMux t3459 (
    .I(seg_21_10_neigh_op_bnl_5_76554),
    .O(seg_21_10_local_g3_5_83972)
  );
  CascadeMux t346 (
    .I(net_54725),
    .O(net_54725_cascademuxed)
  );
  LocalMux t3460 (
    .I(seg_18_10_sp4_h_r_19_69352),
    .O(seg_18_10_local_g0_3_73084)
  );
  Span4Mux_h4 t3461 (
    .I(seg_21_10_sp4_v_b_6_79856),
    .O(seg_18_10_sp4_h_r_19_69352)
  );
  LocalMux t3462 (
    .I(seg_20_9_sp4_r_v_b_33_79980),
    .O(seg_20_9_local_g0_2_79991)
  );
  LocalMux t3463 (
    .I(seg_20_7_sp4_v_b_26_76402),
    .O(seg_20_7_local_g2_2_79761)
  );
  LocalMux t3464 (
    .I(seg_20_9_neigh_op_top_0_76651),
    .O(seg_20_9_local_g1_0_79997)
  );
  LocalMux t3465 (
    .I(seg_20_10_lutff_0_out_76651),
    .O(seg_20_10_local_g3_0_80136)
  );
  LocalMux t3466 (
    .I(seg_21_10_neigh_op_lft_0_76651),
    .O(seg_21_10_local_g0_0_83943)
  );
  LocalMux t3467 (
    .I(seg_20_9_neigh_op_top_3_76654),
    .O(seg_20_9_local_g1_3_80000)
  );
  LocalMux t3468 (
    .I(seg_20_10_lutff_3_out_76654),
    .O(seg_20_10_local_g1_3_80123)
  );
  LocalMux t3469 (
    .I(seg_21_10_neigh_op_lft_3_76654),
    .O(seg_21_10_local_g0_3_83946)
  );
  CascadeMux t347 (
    .I(net_54731),
    .O(net_54731_cascademuxed)
  );
  LocalMux t3470 (
    .I(seg_20_10_lutff_7_out_76658),
    .O(seg_20_10_local_g0_7_80119)
  );
  LocalMux t3471 (
    .I(seg_20_17_sp12_v_b_1_79589),
    .O(seg_20_17_local_g2_1_80990)
  );
  LocalMux t3472 (
    .I(seg_20_10_sp4_v_b_5_76505),
    .O(seg_20_10_local_g1_5_80125)
  );
  Span4Mux_v4 t3473 (
    .I(seg_20_10_sp4_h_r_0_80206),
    .O(seg_20_10_sp4_v_b_5_76505)
  );
  LocalMux t3474 (
    .I(seg_21_10_sp4_h_r_13_80206),
    .O(seg_21_10_local_g1_5_83956)
  );
  LocalMux t3475 (
    .I(seg_20_10_sp4_h_r_10_80208),
    .O(seg_20_10_local_g0_2_80114)
  );
  LocalMux t3476 (
    .I(seg_15_10_sp4_h_r_6_61690),
    .O(seg_15_10_local_g1_6_61602)
  );
  Span4Mux_h4 t3477 (
    .I(seg_19_10_sp4_h_r_3_76800),
    .O(seg_15_10_sp4_h_r_6_61690)
  );
  LocalMux t3478 (
    .I(seg_20_14_sp4_r_v_b_16_80468),
    .O(seg_20_14_local_g3_0_80628)
  );
  Span4Mux_v4 t3479 (
    .I(seg_21_11_sp4_v_b_2_79975),
    .O(seg_20_14_sp4_r_v_b_16_80468)
  );
  CascadeMux t348 (
    .I(net_54737),
    .O(net_54737_cascademuxed)
  );
  LocalMux t3480 (
    .I(seg_20_18_sp4_r_v_b_16_80960),
    .O(seg_20_18_local_g3_0_81120)
  );
  Span4Mux_v4 t3481 (
    .I(seg_21_15_sp4_v_b_5_80468),
    .O(seg_20_18_sp4_r_v_b_16_80960)
  );
  Span4Mux_v4 t3482 (
    .I(seg_21_11_sp4_v_b_2_79975),
    .O(seg_21_15_sp4_v_b_5_80468)
  );
  LocalMux t3483 (
    .I(seg_21_18_sp4_v_b_21_80965),
    .O(seg_21_18_local_g1_5_84940)
  );
  Span4Mux_v4 t3484 (
    .I(seg_21_15_sp4_v_b_5_80468),
    .O(seg_21_18_sp4_v_b_21_80965)
  );
  LocalMux t3485 (
    .I(seg_21_15_sp4_v_b_23_80598),
    .O(seg_21_15_local_g1_7_84573)
  );
  Span4Mux_v4 t3486 (
    .I(seg_21_12_sp4_v_b_7_80101),
    .O(seg_21_15_sp4_v_b_23_80598)
  );
  LocalMux t3487 (
    .I(seg_21_12_sp4_v_b_23_80229),
    .O(seg_21_12_local_g1_7_84204)
  );
  LocalMux t3488 (
    .I(seg_21_13_sp4_v_b_10_80229),
    .O(seg_21_13_local_g1_2_84322)
  );
  LocalMux t3489 (
    .I(seg_21_16_sp4_v_b_23_80721),
    .O(seg_21_16_local_g1_7_84696)
  );
  CascadeMux t349 (
    .I(net_54743),
    .O(net_54743_cascademuxed)
  );
  Span4Mux_v4 t3490 (
    .I(seg_21_13_sp4_v_b_10_80229),
    .O(seg_21_16_sp4_v_b_23_80721)
  );
  LocalMux t3491 (
    .I(seg_18_17_sp4_h_r_28_66380),
    .O(seg_18_17_local_g2_4_73962)
  );
  Span4Mux_h4 t3492 (
    .I(seg_20_17_sp4_v_b_11_77225),
    .O(seg_18_17_sp4_h_r_28_66380)
  );
  Span4Mux_v4 t3493 (
    .I(seg_20_13_sp4_v_b_11_76817),
    .O(seg_20_17_sp4_v_b_11_77225)
  );
  LocalMux t3494 (
    .I(seg_20_13_sp4_v_b_11_76817),
    .O(seg_20_13_local_g1_3_80492)
  );
  GlobalMux t3495 (
    .I(seg_12_0_local_g0_3_48895_i3),
    .O(seg_16_17_glb_netwk_5_10)
  );
  gio2CtrlBuf t3496 (
    .I(seg_12_0_local_g0_3_48895_i2),
    .O(seg_12_0_local_g0_3_48895_i3)
  );
  ICE_GB t3497 (
    .GLOBALBUFFEROUTPUT(seg_12_0_local_g0_3_48895_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_12_0_local_g0_3_48895_i1)
  );
  IoInMux t3498 (
    .I(seg_12_0_local_g0_3_48895),
    .O(seg_12_0_local_g0_3_48895_i1)
  );
  LocalMux t3499 (
    .I(seg_12_0_span4_vert_19_45240),
    .O(seg_12_0_local_g0_3_48895)
  );
  CascadeMux t35 (
    .I(net_20982),
    .O(net_20982_cascademuxed)
  );
  CascadeMux t350 (
    .I(net_54824),
    .O(net_54824_cascademuxed)
  );
  Span4Mux_v4 t3500 (
    .I(seg_12_2_sp4_h_r_6_49215),
    .O(seg_12_0_span4_vert_19_45240)
  );
  Span4Mux_h4 t3501 (
    .I(seg_16_2_sp4_h_r_6_64537),
    .O(seg_12_2_sp4_h_r_6_49215)
  );
  Span4Mux_h4 t3502 (
    .I(seg_20_2_sp4_v_t_43_76100),
    .O(seg_16_2_sp4_h_r_6_64537)
  );
  Span4Mux_v4 t3503 (
    .I(seg_20_6_sp4_v_t_43_76508),
    .O(seg_20_2_sp4_v_t_43_76100)
  );
  LocalMux t3504 (
    .I(seg_20_12_neigh_op_bot_5_76758),
    .O(seg_20_12_local_g1_5_80371)
  );
  LocalMux t3505 (
    .I(seg_21_12_neigh_op_lft_0_76855),
    .O(seg_21_12_local_g0_0_84189)
  );
  LocalMux t3506 (
    .I(seg_20_12_lutff_1_out_76856),
    .O(seg_20_12_local_g2_1_80375)
  );
  LocalMux t3507 (
    .I(seg_20_12_lutff_2_out_76857),
    .O(seg_20_12_local_g1_2_80368)
  );
  LocalMux t3508 (
    .I(seg_20_12_lutff_3_out_76858),
    .O(seg_20_12_local_g1_3_80369)
  );
  LocalMux t3509 (
    .I(seg_20_13_neigh_op_bot_4_76859),
    .O(seg_20_13_local_g1_4_80493)
  );
  CascadeMux t351 (
    .I(net_54830),
    .O(net_54830_cascademuxed)
  );
  LocalMux t3510 (
    .I(seg_20_12_lutff_5_out_76860),
    .O(seg_20_12_local_g2_5_80379)
  );
  LocalMux t3511 (
    .I(seg_20_12_lutff_6_out_76861),
    .O(seg_20_12_local_g3_6_80388)
  );
  LocalMux t3512 (
    .I(seg_21_12_neigh_op_lft_7_76862),
    .O(seg_21_12_local_g0_7_84196)
  );
  LocalMux t3513 (
    .I(seg_21_14_neigh_op_bnl_0_76957),
    .O(seg_21_14_local_g3_0_84459)
  );
  LocalMux t3514 (
    .I(seg_21_13_neigh_op_lft_4_76961),
    .O(seg_21_13_local_g1_4_84324)
  );
  LocalMux t3515 (
    .I(seg_20_14_neigh_op_bot_7_76964),
    .O(seg_20_14_local_g1_7_80619)
  );
  LocalMux t3516 (
    .I(seg_18_13_sp4_h_r_10_73546),
    .O(seg_18_13_local_g0_2_73452)
  );
  LocalMux t3517 (
    .I(seg_18_13_sp4_h_r_12_69714),
    .O(seg_18_13_local_g1_4_73462)
  );
  LocalMux t3518 (
    .I(seg_21_15_sp4_v_b_31_80716),
    .O(seg_21_15_local_g3_7_84589)
  );
  Span4Mux_v4 t3519 (
    .I(seg_21_13_sp4_h_l_42_69722),
    .O(seg_21_15_sp4_v_b_31_80716)
  );
  CascadeMux t352 (
    .I(net_54836),
    .O(net_54836_cascademuxed)
  );
  LocalMux t3520 (
    .I(seg_18_14_sp4_h_r_35_66008),
    .O(seg_18_14_local_g2_3_73592)
  );
  Span4Mux_h4 t3521 (
    .I(seg_20_14_sp4_v_b_11_76919),
    .O(seg_18_14_sp4_h_r_35_66008)
  );
  LocalMux t3522 (
    .I(seg_20_15_sp4_v_b_4_77016),
    .O(seg_20_15_local_g1_4_80739)
  );
  LocalMux t3523 (
    .I(seg_20_14_lutff_0_out_77059),
    .O(seg_20_14_local_g1_0_80612)
  );
  LocalMux t3524 (
    .I(seg_20_13_neigh_op_top_1_77060),
    .O(seg_20_13_local_g0_1_80482)
  );
  LocalMux t3525 (
    .I(seg_20_13_neigh_op_top_2_77061),
    .O(seg_20_13_local_g0_2_80483)
  );
  LocalMux t3526 (
    .I(seg_21_14_neigh_op_lft_3_77062),
    .O(seg_21_14_local_g0_3_84438)
  );
  LocalMux t3527 (
    .I(seg_20_13_neigh_op_top_4_77063),
    .O(seg_20_13_local_g0_4_80485)
  );
  LocalMux t3528 (
    .I(seg_20_14_lutff_5_out_77064),
    .O(seg_20_14_local_g0_5_80609)
  );
  LocalMux t3529 (
    .I(seg_20_13_neigh_op_top_6_77065),
    .O(seg_20_13_local_g1_6_80495)
  );
  CascadeMux t353 (
    .I(net_54842),
    .O(net_54842_cascademuxed)
  );
  LocalMux t3530 (
    .I(seg_21_14_neigh_op_lft_7_77066),
    .O(seg_21_14_local_g0_7_84442)
  );
  LocalMux t3531 (
    .I(seg_21_15_neigh_op_lft_0_77161),
    .O(seg_21_15_local_g1_0_84566)
  );
  LocalMux t3532 (
    .I(seg_20_14_neigh_op_top_1_77162),
    .O(seg_20_14_local_g1_1_80613)
  );
  LocalMux t3533 (
    .I(seg_21_15_neigh_op_lft_2_77163),
    .O(seg_21_15_local_g1_2_84568)
  );
  LocalMux t3534 (
    .I(seg_21_15_neigh_op_lft_3_77164),
    .O(seg_21_15_local_g0_3_84561)
  );
  LocalMux t3535 (
    .I(seg_20_15_lutff_4_out_77165),
    .O(seg_20_15_local_g0_4_80731)
  );
  LocalMux t3536 (
    .I(seg_21_15_neigh_op_lft_5_77166),
    .O(seg_21_15_local_g0_5_84563)
  );
  LocalMux t3537 (
    .I(seg_20_12_sp4_h_r_6_80460),
    .O(seg_20_12_local_g1_6_80372)
  );
  Span4Mux_h4 t3538 (
    .I(seg_20_12_sp4_v_t_36_77113),
    .O(seg_20_12_sp4_h_r_6_80460)
  );
  LocalMux t3539 (
    .I(seg_20_14_sp4_v_b_27_77115),
    .O(seg_20_14_local_g2_3_80623)
  );
  CascadeMux t354 (
    .I(net_54848),
    .O(net_54848_cascademuxed)
  );
  LocalMux t3540 (
    .I(seg_19_16_neigh_op_rgt_1_77264),
    .O(seg_19_16_local_g3_1_77358)
  );
  LocalMux t3541 (
    .I(seg_20_16_lutff_1_out_77264),
    .O(seg_20_16_local_g1_1_80859)
  );
  LocalMux t3542 (
    .I(seg_21_17_neigh_op_bnl_1_77264),
    .O(seg_21_17_local_g3_1_84829)
  );
  LocalMux t3543 (
    .I(seg_19_16_neigh_op_rgt_2_77265),
    .O(seg_19_16_local_g3_2_77359)
  );
  LocalMux t3544 (
    .I(seg_20_16_lutff_2_out_77265),
    .O(seg_20_16_local_g2_2_80868)
  );
  LocalMux t3545 (
    .I(seg_21_17_neigh_op_bnl_2_77265),
    .O(seg_21_17_local_g3_2_84830)
  );
  LocalMux t3546 (
    .I(seg_19_16_neigh_op_rgt_3_77266),
    .O(seg_19_16_local_g3_3_77360)
  );
  LocalMux t3547 (
    .I(seg_20_16_lutff_3_out_77266),
    .O(seg_20_16_local_g3_3_80877)
  );
  LocalMux t3548 (
    .I(seg_21_17_neigh_op_bnl_3_77266),
    .O(seg_21_17_local_g3_3_84831)
  );
  LocalMux t3549 (
    .I(seg_19_16_neigh_op_rgt_4_77267),
    .O(seg_19_16_local_g3_4_77361)
  );
  CascadeMux t355 (
    .I(net_54854),
    .O(net_54854_cascademuxed)
  );
  LocalMux t3550 (
    .I(seg_20_16_lutff_4_out_77267),
    .O(seg_20_16_local_g1_4_80862)
  );
  LocalMux t3551 (
    .I(seg_20_17_neigh_op_bot_4_77267),
    .O(seg_20_17_local_g0_4_80977)
  );
  LocalMux t3552 (
    .I(seg_19_16_neigh_op_rgt_5_77268),
    .O(seg_19_16_local_g3_5_77362)
  );
  LocalMux t3553 (
    .I(seg_20_16_lutff_5_out_77268),
    .O(seg_20_16_local_g2_5_80871)
  );
  LocalMux t3554 (
    .I(seg_20_17_neigh_op_bot_5_77268),
    .O(seg_20_17_local_g0_5_80978)
  );
  LocalMux t3555 (
    .I(seg_19_16_neigh_op_rgt_6_77269),
    .O(seg_19_16_local_g3_6_77363)
  );
  LocalMux t3556 (
    .I(seg_20_16_lutff_6_out_77269),
    .O(seg_20_16_local_g1_6_80864)
  );
  LocalMux t3557 (
    .I(seg_21_17_neigh_op_bnl_6_77269),
    .O(seg_21_17_local_g3_6_84834)
  );
  LocalMux t3558 (
    .I(seg_19_16_neigh_op_rgt_7_77270),
    .O(seg_19_16_local_g3_7_77364)
  );
  LocalMux t3559 (
    .I(seg_20_16_lutff_7_out_77270),
    .O(seg_20_16_local_g3_7_80881)
  );
  CascadeMux t356 (
    .I(net_54860),
    .O(net_54860_cascademuxed)
  );
  LocalMux t3560 (
    .I(seg_21_17_neigh_op_bnl_7_77270),
    .O(seg_21_17_local_g2_7_84827)
  );
  LocalMux t3561 (
    .I(seg_19_18_sp4_r_v_b_34_77532),
    .O(seg_19_18_local_g0_1_77538)
  );
  Span4Mux_v4 t3562 (
    .I(seg_20_16_sp4_h_r_4_80950),
    .O(seg_19_18_sp4_r_v_b_34_77532)
  );
  LocalMux t3563 (
    .I(seg_19_18_sp4_h_r_32_70338),
    .O(seg_19_18_local_g2_0_77553)
  );
  Span4Mux_h4 t3564 (
    .I(seg_21_18_sp4_v_b_3_80835),
    .O(seg_19_18_sp4_h_r_32_70338)
  );
  LocalMux t3565 (
    .I(seg_19_18_sp4_h_r_31_70337),
    .O(seg_19_18_local_g3_7_77568)
  );
  Span4Mux_h4 t3566 (
    .I(seg_21_18_sp4_v_b_7_80839),
    .O(seg_19_18_sp4_h_r_31_70337)
  );
  LocalMux t3567 (
    .I(seg_19_14_sp4_r_v_b_34_77124),
    .O(seg_19_14_local_g2_2_77147)
  );
  LocalMux t3568 (
    .I(seg_19_14_sp4_r_v_b_38_77217),
    .O(seg_19_14_local_g2_6_77151)
  );
  LocalMux t3569 (
    .I(seg_19_14_sp4_r_v_b_26_77116),
    .O(seg_19_14_local_g0_2_77131)
  );
  CascadeMux t357 (
    .I(net_54866),
    .O(net_54866_cascademuxed)
  );
  LocalMux t3570 (
    .I(seg_19_14_sp4_r_v_b_44_77223),
    .O(seg_19_14_local_g3_4_77157)
  );
  LocalMux t3571 (
    .I(seg_19_14_sp4_r_v_b_0_76910),
    .O(seg_19_14_local_g1_0_77137)
  );
  Span4Mux_v4 t3572 (
    .I(seg_20_14_sp4_v_t_41_77322),
    .O(seg_19_14_sp4_r_v_b_0_76910)
  );
  LocalMux t3573 (
    .I(seg_19_18_sp4_r_v_b_4_77322),
    .O(seg_19_18_local_g1_4_77549)
  );
  LocalMux t3574 (
    .I(seg_19_18_sp4_r_v_b_10_77328),
    .O(seg_19_18_local_g2_2_77555)
  );
  LocalMux t3575 (
    .I(seg_19_18_sp4_r_v_b_14_77421),
    .O(seg_19_18_local_g2_6_77559)
  );
  LocalMux t3576 (
    .I(seg_19_18_sp4_r_v_b_16_77423),
    .O(seg_19_18_local_g3_0_77561)
  );
  LocalMux t3577 (
    .I(seg_19_14_sp4_r_v_b_30_77120),
    .O(seg_19_14_local_g0_6_77135)
  );
  LocalMux t3578 (
    .I(seg_19_14_sp4_r_v_b_32_77122),
    .O(seg_19_14_local_g0_3_77132)
  );
  LocalMux t3579 (
    .I(seg_21_16_neigh_op_tnl_1_77366),
    .O(seg_21_16_local_g3_1_84706)
  );
  CascadeMux t358 (
    .I(net_55076),
    .O(net_55076_cascademuxed)
  );
  LocalMux t3580 (
    .I(seg_21_17_neigh_op_lft_2_77367),
    .O(seg_21_17_local_g1_2_84814)
  );
  LocalMux t3581 (
    .I(seg_20_17_lutff_3_out_77368),
    .O(seg_20_17_local_g2_3_80992)
  );
  LocalMux t3582 (
    .I(seg_20_17_lutff_5_out_77370),
    .O(seg_20_17_local_g3_5_81002)
  );
  LocalMux t3583 (
    .I(seg_20_17_lutff_6_out_77371),
    .O(seg_20_17_local_g0_6_80979)
  );
  LocalMux t3584 (
    .I(seg_20_17_lutff_7_out_77372),
    .O(seg_20_17_local_g0_7_80980)
  );
  LocalMux t3585 (
    .I(seg_21_14_sp4_v_b_36_80710),
    .O(seg_21_14_local_g3_4_84463)
  );
  LocalMux t3586 (
    .I(seg_21_14_sp4_v_b_44_80718),
    .O(seg_21_14_local_g2_4_84455)
  );
  LocalMux t3587 (
    .I(seg_21_18_neigh_op_lft_1_77468),
    .O(seg_21_18_local_g0_1_84928)
  );
  LocalMux t3588 (
    .I(seg_21_18_neigh_op_lft_3_77470),
    .O(seg_21_18_local_g1_3_84938)
  );
  LocalMux t3589 (
    .I(seg_21_18_neigh_op_lft_4_77471),
    .O(seg_21_18_local_g1_4_84939)
  );
  CascadeMux t359 (
    .I(net_55082),
    .O(net_55082_cascademuxed)
  );
  LocalMux t3590 (
    .I(seg_20_18_lutff_7_out_77474),
    .O(seg_20_18_local_g2_7_81119)
  );
  LocalMux t3591 (
    .I(seg_21_14_sp4_v_b_30_80594),
    .O(seg_21_14_local_g3_6_84465)
  );
  Span4Mux_v4 t3592 (
    .I(seg_21_16_sp4_v_t_38_81081),
    .O(seg_21_14_sp4_v_b_30_80594)
  );
  LocalMux t3593 (
    .I(seg_20_18_neigh_op_top_6_77575),
    .O(seg_20_18_local_g1_6_81110)
  );
  LocalMux t3594 (
    .I(seg_20_18_neigh_op_top_7_77576),
    .O(seg_20_18_local_g1_7_81111)
  );
  LocalMux t3595 (
    .I(seg_20_6_neigh_op_rgt_5_79584),
    .O(seg_20_6_local_g3_5_79649)
  );
  LocalMux t3596 (
    .I(seg_20_7_neigh_op_bnr_5_79584),
    .O(seg_20_7_local_g1_5_79756)
  );
  LocalMux t3597 (
    .I(seg_21_9_sp12_v_b_5_82776),
    .O(seg_21_9_local_g3_5_83849)
  );
  LocalMux t3598 (
    .I(seg_21_14_sp4_v_b_4_80346),
    .O(seg_21_14_local_g0_4_84439)
  );
  Span4Mux_v4 t3599 (
    .I(seg_21_10_sp4_v_b_4_79854),
    .O(seg_21_14_sp4_v_b_4_80346)
  );
  CascadeMux t36 (
    .I(net_21099),
    .O(net_21099_cascademuxed)
  );
  CascadeMux t360 (
    .I(net_55094),
    .O(net_55094_cascademuxed)
  );
  Span4Mux_v4 t3600 (
    .I(seg_21_6_sp4_h_r_10_83547),
    .O(seg_21_10_sp4_v_b_4_79854)
  );
  LocalMux t3601 (
    .I(seg_17_6_sp4_h_r_29_61197),
    .O(seg_17_6_local_g3_5_68787)
  );
  Span4Mux_h4 t3602 (
    .I(seg_19_6_sp4_h_r_2_76391),
    .O(seg_17_6_sp4_h_r_29_61197)
  );
  LocalMux t3603 (
    .I(seg_17_5_sp4_r_v_b_12_68495),
    .O(seg_17_5_local_g2_4_68655)
  );
  Span4Mux_v4 t3604 (
    .I(seg_18_6_sp4_h_l_42_57369),
    .O(seg_17_5_sp4_r_v_b_12_68495)
  );
  Span4Mux_h4 t3605 (
    .I(seg_18_6_sp4_h_r_7_72692),
    .O(seg_18_6_sp4_h_l_42_57369)
  );
  LocalMux t3606 (
    .I(seg_18_5_sp4_v_b_13_68496),
    .O(seg_18_5_local_g1_5_72479)
  );
  Span4Mux_v4 t3607 (
    .I(seg_18_6_sp4_h_r_7_72692),
    .O(seg_18_5_sp4_v_b_13_68496)
  );
  LocalMux t3608 (
    .I(seg_18_6_sp4_h_r_7_72692),
    .O(seg_18_6_local_g0_7_72596)
  );
  LocalMux t3609 (
    .I(seg_18_6_sp4_h_r_4_72689),
    .O(seg_18_6_local_g0_4_72593)
  );
  CascadeMux t361 (
    .I(net_55106),
    .O(net_55106_cascademuxed)
  );
  Span4Mux_h4 t3610 (
    .I(seg_22_6_sp4_v_b_11_83198),
    .O(seg_18_6_sp4_h_r_4_72689)
  );
  LocalMux t3611 (
    .I(seg_23_9_sp4_h_r_13_87745),
    .O(seg_23_9_local_g1_5_91495)
  );
  Span4Mux_h4 t3612 (
    .I(seg_22_9_sp4_v_b_6_83564),
    .O(seg_23_9_sp4_h_r_13_87745)
  );
  LocalMux t3613 (
    .I(seg_22_0_span4_vert_18_82916),
    .O(seg_22_0_local_g1_2_86579)
  );
  Span4Mux_v4 t3614 (
    .I(seg_22_2_sp4_v_t_42_83194),
    .O(seg_22_0_span4_vert_18_82916)
  );
  LocalMux t3615 (
    .I(seg_21_14_sp4_v_b_9_80349),
    .O(seg_21_14_local_g0_1_84436)
  );
  Span4Mux_v4 t3616 (
    .I(seg_21_10_sp4_v_b_1_79849),
    .O(seg_21_14_sp4_v_b_9_80349)
  );
  Span4Mux_v4 t3617 (
    .I(seg_21_6_sp4_v_b_10_79368),
    .O(seg_21_10_sp4_v_b_1_79849)
  );
  LocalMux t3618 (
    .I(seg_20_9_sp4_r_v_b_7_79732),
    .O(seg_20_9_local_g1_7_80004)
  );
  LocalMux t3619 (
    .I(seg_22_9_sp4_h_r_12_83915),
    .O(seg_22_9_local_g0_4_87655)
  );
  CascadeMux t362 (
    .I(net_55112),
    .O(net_55112_cascademuxed)
  );
  Span4Mux_h4 t3620 (
    .I(seg_21_9_sp4_v_b_7_79732),
    .O(seg_22_9_sp4_h_r_12_83915)
  );
  LocalMux t3621 (
    .I(seg_21_9_lutff_0_out_79948),
    .O(seg_21_9_local_g1_0_83828)
  );
  LocalMux t3622 (
    .I(seg_21_9_lutff_2_out_79950),
    .O(seg_21_9_local_g0_2_83822)
  );
  LocalMux t3623 (
    .I(seg_21_14_sp12_v_b_11_83667),
    .O(seg_21_14_local_g3_3_84462)
  );
  LocalMux t3624 (
    .I(seg_23_9_sp4_h_r_24_83914),
    .O(seg_23_9_local_g3_0_91506)
  );
  LocalMux t3625 (
    .I(seg_23_9_sp4_r_v_b_3_91221),
    .O(seg_23_9_local_g1_3_91493)
  );
  Span4Mux_v4 t3626 (
    .I(seg_24_9_sp4_h_l_44_80094),
    .O(seg_23_9_sp4_r_v_b_3_91221)
  );
  LocalMux t3627 (
    .I(seg_22_9_sp4_r_v_b_10_87399),
    .O(seg_22_9_local_g2_2_87669)
  );
  Span4Mux_v4 t3628 (
    .I(seg_23_9_sp4_h_l_41_76699),
    .O(seg_22_9_sp4_r_v_b_10_87399)
  );
  LocalMux t3629 (
    .I(seg_21_15_sp4_v_b_18_80593),
    .O(seg_21_15_local_g0_2_84560)
  );
  CascadeMux t363 (
    .I(net_55217),
    .O(net_55217_cascademuxed)
  );
  Span4Mux_v4 t3630 (
    .I(seg_21_12_sp4_h_r_7_84292),
    .O(seg_21_15_sp4_v_b_18_80593)
  );
  Span4Mux_h4 t3631 (
    .I(seg_21_12_sp4_v_b_1_80095),
    .O(seg_21_12_sp4_h_r_7_84292)
  );
  LocalMux t3632 (
    .I(seg_21_10_lutff_0_out_80071),
    .O(seg_21_10_local_g3_0_83967)
  );
  LocalMux t3633 (
    .I(seg_20_10_neigh_op_rgt_1_80072),
    .O(seg_20_10_local_g3_1_80137)
  );
  LocalMux t3634 (
    .I(seg_20_10_neigh_op_rgt_4_80075),
    .O(seg_20_10_local_g2_4_80132)
  );
  LocalMux t3635 (
    .I(seg_20_10_neigh_op_rgt_4_80075),
    .O(seg_20_10_local_g3_4_80140)
  );
  LocalMux t3636 (
    .I(seg_21_10_lutff_4_out_80075),
    .O(seg_21_10_local_g2_4_83963)
  );
  LocalMux t3637 (
    .I(seg_21_18_sp12_v_b_2_83666),
    .O(seg_21_18_local_g3_2_84953)
  );
  LocalMux t3638 (
    .I(seg_21_10_sp4_h_r_10_84039),
    .O(seg_21_10_local_g0_2_83945)
  );
  LocalMux t3639 (
    .I(seg_20_14_sp4_v_b_1_76909),
    .O(seg_20_14_local_g0_1_80605)
  );
  CascadeMux t364 (
    .I(net_55223),
    .O(net_55223_cascademuxed)
  );
  Span4Mux_v4 t3640 (
    .I(seg_20_10_sp4_h_r_7_80215),
    .O(seg_20_14_sp4_v_b_1_76909)
  );
  LocalMux t3641 (
    .I(seg_17_17_sp4_v_b_12_66140),
    .O(seg_17_17_local_g1_4_70123)
  );
  Span4Mux_v4 t3642 (
    .I(seg_17_14_sp4_v_b_10_65659),
    .O(seg_17_17_sp4_v_b_12_66140)
  );
  Span4Mux_v4 t3643 (
    .I(seg_17_10_sp4_h_r_10_69346),
    .O(seg_17_14_sp4_v_b_10_65659)
  );
  Span4Mux_h4 t3644 (
    .I(seg_21_10_sp4_h_r_2_84041),
    .O(seg_17_10_sp4_h_r_10_69346)
  );
  LocalMux t3645 (
    .I(seg_20_17_sp4_r_v_b_15_80836),
    .O(seg_20_17_local_g2_7_80996)
  );
  Span4Mux_v4 t3646 (
    .I(seg_21_14_sp4_v_b_2_80344),
    .O(seg_20_17_sp4_r_v_b_15_80836)
  );
  Span4Mux_v4 t3647 (
    .I(seg_21_10_sp4_h_r_2_84041),
    .O(seg_21_14_sp4_v_b_2_80344)
  );
  LocalMux t3648 (
    .I(seg_21_13_sp4_v_b_15_80344),
    .O(seg_21_13_local_g0_7_84319)
  );
  Span4Mux_v4 t3649 (
    .I(seg_21_10_sp4_h_r_2_84041),
    .O(seg_21_13_sp4_v_b_15_80344)
  );
  CascadeMux t365 (
    .I(net_55229),
    .O(net_55229_cascademuxed)
  );
  LocalMux t3650 (
    .I(seg_15_10_sp4_h_r_0_61682),
    .O(seg_15_10_local_g0_0_61588)
  );
  Span4Mux_h4 t3651 (
    .I(seg_19_10_sp4_h_r_0_76795),
    .O(seg_15_10_sp4_h_r_0_61682)
  );
  LocalMux t3652 (
    .I(seg_18_17_sp4_r_v_b_20_73810),
    .O(seg_18_17_local_g3_4_73970)
  );
  Span4Mux_v4 t3653 (
    .I(seg_19_14_sp4_v_b_6_73317),
    .O(seg_18_17_sp4_r_v_b_20_73810)
  );
  Span4Mux_v4 t3654 (
    .I(seg_19_10_sp4_h_r_0_76795),
    .O(seg_19_14_sp4_v_b_6_73317)
  );
  LocalMux t3655 (
    .I(seg_15_10_sp4_h_r_10_61684),
    .O(seg_15_10_local_g1_2_61598)
  );
  Span4Mux_h4 t3656 (
    .I(seg_19_10_sp4_h_r_10_76797),
    .O(seg_15_10_sp4_h_r_10_61684)
  );
  LocalMux t3657 (
    .I(seg_18_13_sp4_r_v_b_17_73315),
    .O(seg_18_13_local_g3_1_73475)
  );
  Span4Mux_v4 t3658 (
    .I(seg_19_10_sp4_h_r_10_76797),
    .O(seg_18_13_sp4_r_v_b_17_73315)
  );
  LocalMux t3659 (
    .I(seg_18_14_sp4_r_v_b_10_73321),
    .O(seg_18_14_local_g2_2_73591)
  );
  CascadeMux t366 (
    .I(net_55235),
    .O(net_55235_cascademuxed)
  );
  Span4Mux_v4 t3660 (
    .I(seg_19_10_sp4_h_r_10_76797),
    .O(seg_18_14_sp4_r_v_b_10_73321)
  );
  LocalMux t3661 (
    .I(seg_18_18_sp4_r_v_b_10_73813),
    .O(seg_18_18_local_g2_2_74083)
  );
  Span4Mux_v4 t3662 (
    .I(seg_19_14_sp4_v_b_10_73321),
    .O(seg_18_18_sp4_r_v_b_10_73813)
  );
  Span4Mux_v4 t3663 (
    .I(seg_19_10_sp4_h_r_10_76797),
    .O(seg_19_14_sp4_v_b_10_73321)
  );
  LocalMux t3664 (
    .I(seg_20_18_sp4_r_v_b_8_80842),
    .O(seg_20_18_local_g2_0_81112)
  );
  Span4Mux_v4 t3665 (
    .I(seg_21_14_sp4_v_b_8_80350),
    .O(seg_20_18_sp4_r_v_b_8_80842)
  );
  Span4Mux_v4 t3666 (
    .I(seg_21_10_sp4_h_r_8_84047),
    .O(seg_21_14_sp4_v_b_8_80350)
  );
  LocalMux t3667 (
    .I(seg_21_18_sp4_v_b_8_80842),
    .O(seg_21_18_local_g1_0_84935)
  );
  Span4Mux_v4 t3668 (
    .I(seg_21_14_sp4_v_b_8_80350),
    .O(seg_21_18_sp4_v_b_8_80842)
  );
  LocalMux t3669 (
    .I(seg_21_15_sp4_r_v_b_12_84418),
    .O(seg_21_15_local_g2_4_84578)
  );
  CascadeMux t367 (
    .I(net_55457),
    .O(net_55457_cascademuxed)
  );
  Span4Mux_v4 t3670 (
    .I(seg_22_12_sp4_v_b_1_83926),
    .O(seg_21_15_sp4_r_v_b_12_84418)
  );
  LocalMux t3671 (
    .I(seg_20_15_sp4_r_v_b_10_80475),
    .O(seg_20_15_local_g2_2_80745)
  );
  Span4Mux_v4 t3672 (
    .I(seg_21_11_sp4_v_b_7_79978),
    .O(seg_20_15_sp4_r_v_b_10_80475)
  );
  LocalMux t3673 (
    .I(seg_20_14_sp4_r_v_b_24_80588),
    .O(seg_20_14_local_g0_0_80604)
  );
  Span4Mux_v4 t3674 (
    .I(seg_21_12_sp4_v_b_0_80096),
    .O(seg_20_14_sp4_r_v_b_24_80588)
  );
  LocalMux t3675 (
    .I(seg_17_15_sp4_v_b_14_65896),
    .O(seg_17_15_local_g1_6_69879)
  );
  Span4Mux_v4 t3676 (
    .I(seg_17_12_sp4_h_r_3_69595),
    .O(seg_17_15_sp4_v_b_14_65896)
  );
  Span4Mux_h4 t3677 (
    .I(seg_21_12_sp4_v_b_10_80106),
    .O(seg_17_12_sp4_h_r_3_69595)
  );
  LocalMux t3678 (
    .I(seg_20_12_sp4_r_v_b_10_80106),
    .O(seg_20_12_local_g2_2_80376)
  );
  LocalMux t3679 (
    .I(seg_21_15_sp4_v_b_12_80587),
    .O(seg_21_15_local_g0_4_84562)
  );
  CascadeMux t368 (
    .I(net_55481),
    .O(net_55481_cascademuxed)
  );
  Span4Mux_v4 t3680 (
    .I(seg_21_12_sp4_v_b_10_80106),
    .O(seg_21_15_sp4_v_b_12_80587)
  );
  LocalMux t3681 (
    .I(seg_21_16_sp4_v_b_1_80587),
    .O(seg_21_16_local_g0_1_84682)
  );
  Span4Mux_v4 t3682 (
    .I(seg_21_12_sp4_v_b_10_80106),
    .O(seg_21_16_sp4_v_b_1_80587)
  );
  LocalMux t3683 (
    .I(seg_20_13_sp4_r_v_b_5_80222),
    .O(seg_20_13_local_g1_5_80494)
  );
  LocalMux t3684 (
    .I(seg_20_17_sp4_r_v_b_5_80714),
    .O(seg_20_17_local_g1_5_80986)
  );
  Span4Mux_v4 t3685 (
    .I(seg_21_13_sp4_v_b_5_80222),
    .O(seg_20_17_sp4_r_v_b_5_80714)
  );
  LocalMux t3686 (
    .I(seg_21_12_sp4_v_b_16_80222),
    .O(seg_21_12_local_g1_0_84197)
  );
  LocalMux t3687 (
    .I(seg_21_13_sp4_v_b_5_80222),
    .O(seg_21_13_local_g1_5_84325)
  );
  LocalMux t3688 (
    .I(seg_21_15_sp4_v_b_32_80719),
    .O(seg_21_15_local_g3_0_84582)
  );
  Span4Mux_v4 t3689 (
    .I(seg_21_13_sp4_v_b_5_80222),
    .O(seg_21_15_sp4_v_b_32_80719)
  );
  CascadeMux t369 (
    .I(net_56066),
    .O(net_56066_cascademuxed)
  );
  LocalMux t3690 (
    .I(seg_21_13_neigh_op_bot_2_80319),
    .O(seg_21_13_local_g0_2_84314)
  );
  LocalMux t3691 (
    .I(seg_20_12_neigh_op_rgt_7_80324),
    .O(seg_20_12_local_g3_7_80389)
  );
  LocalMux t3692 (
    .I(seg_21_14_sp4_v_b_18_80470),
    .O(seg_21_14_local_g0_2_84437)
  );
  LocalMux t3693 (
    .I(seg_21_13_lutff_1_out_80441),
    .O(seg_21_13_local_g1_1_84321)
  );
  LocalMux t3694 (
    .I(seg_21_14_neigh_op_bot_2_80442),
    .O(seg_21_14_local_g1_2_84445)
  );
  LocalMux t3695 (
    .I(seg_21_13_lutff_6_out_80446),
    .O(seg_21_13_local_g2_6_84334)
  );
  LocalMux t3696 (
    .I(seg_20_14_neigh_op_bnr_7_80447),
    .O(seg_20_14_local_g0_7_80611)
  );
  LocalMux t3697 (
    .I(seg_21_15_sp4_r_v_b_17_84423),
    .O(seg_21_15_local_g3_1_84583)
  );
  LocalMux t3698 (
    .I(seg_21_15_sp4_v_b_8_80473),
    .O(seg_21_15_local_g0_0_84558)
  );
  LocalMux t3699 (
    .I(seg_21_15_sp4_v_b_14_80589),
    .O(seg_21_15_local_g1_6_84572)
  );
  CascadeMux t37 (
    .I(net_21111),
    .O(net_21111_cascademuxed)
  );
  CascadeMux t370 (
    .I(net_56084),
    .O(net_56084_cascademuxed)
  );
  LocalMux t3700 (
    .I(seg_21_14_lutff_1_out_80564),
    .O(seg_21_14_local_g2_1_84452)
  );
  LocalMux t3701 (
    .I(seg_21_14_lutff_2_out_80565),
    .O(seg_21_14_local_g2_2_84453)
  );
  LocalMux t3702 (
    .I(seg_21_14_lutff_3_out_80566),
    .O(seg_21_14_local_g2_3_84454)
  );
  LocalMux t3703 (
    .I(seg_21_14_lutff_4_out_80567),
    .O(seg_21_14_local_g1_4_84447)
  );
  LocalMux t3704 (
    .I(seg_21_14_lutff_5_out_80568),
    .O(seg_21_14_local_g2_5_84456)
  );
  LocalMux t3705 (
    .I(seg_21_14_lutff_7_out_80570),
    .O(seg_21_14_local_g2_7_84458)
  );
  LocalMux t3706 (
    .I(seg_21_6_sp4_v_b_17_79485),
    .O(seg_21_6_local_g1_1_83460)
  );
  Span4Mux_v4 t3707 (
    .I(seg_21_7_sp4_v_t_41_79977),
    .O(seg_21_6_sp4_v_b_17_79485)
  );
  Span4Mux_v4 t3708 (
    .I(seg_21_11_sp4_v_t_36_80464),
    .O(seg_21_7_sp4_v_t_41_79977)
  );
  LocalMux t3709 (
    .I(seg_21_15_sp4_v_b_21_80596),
    .O(seg_21_15_local_g1_5_84571)
  );
  CascadeMux t371 (
    .I(net_56090),
    .O(net_56090_cascademuxed)
  );
  LocalMux t3710 (
    .I(seg_21_14_neigh_op_top_0_80686),
    .O(seg_21_14_local_g1_0_84443)
  );
  LocalMux t3711 (
    .I(seg_21_14_neigh_op_top_1_80687),
    .O(seg_21_14_local_g1_1_84444)
  );
  LocalMux t3712 (
    .I(seg_21_15_lutff_2_out_80688),
    .O(seg_21_15_local_g3_2_84584)
  );
  LocalMux t3713 (
    .I(seg_21_15_lutff_3_out_80689),
    .O(seg_21_15_local_g3_3_84585)
  );
  LocalMux t3714 (
    .I(seg_21_15_lutff_4_out_80690),
    .O(seg_21_15_local_g1_4_84570)
  );
  LocalMux t3715 (
    .I(seg_21_14_neigh_op_top_5_80691),
    .O(seg_21_14_local_g1_5_84448)
  );
  LocalMux t3716 (
    .I(seg_21_15_lutff_6_out_80692),
    .O(seg_21_15_local_g0_6_84564)
  );
  LocalMux t3717 (
    .I(seg_21_14_neigh_op_top_7_80693),
    .O(seg_21_14_local_g1_7_84450)
  );
  LocalMux t3718 (
    .I(seg_21_15_neigh_op_top_3_80812),
    .O(seg_21_15_local_g1_3_84569)
  );
  LocalMux t3719 (
    .I(seg_21_17_neigh_op_bot_4_80813),
    .O(seg_21_17_local_g0_4_84808)
  );
  CascadeMux t372 (
    .I(net_56821),
    .O(net_56821_cascademuxed)
  );
  LocalMux t3720 (
    .I(seg_21_16_lutff_6_out_80815),
    .O(seg_21_16_local_g3_6_84711)
  );
  LocalMux t3721 (
    .I(seg_19_13_sp4_v_b_37_73557),
    .O(seg_19_13_local_g2_5_77048)
  );
  Span4Mux_v4 t3722 (
    .I(seg_19_16_sp4_h_r_0_77407),
    .O(seg_19_13_sp4_v_b_37_73557)
  );
  LocalMux t3723 (
    .I(seg_19_15_sp4_v_b_13_73557),
    .O(seg_19_15_local_g0_5_77236)
  );
  Span4Mux_v4 t3724 (
    .I(seg_19_16_sp4_h_r_0_77407),
    .O(seg_19_15_sp4_v_b_13_73557)
  );
  LocalMux t3725 (
    .I(seg_19_17_sp4_v_b_37_74049),
    .O(seg_19_17_local_g2_5_77456)
  );
  Span4Mux_v4 t3726 (
    .I(seg_19_16_sp4_h_r_0_77407),
    .O(seg_19_17_sp4_v_b_37_74049)
  );
  LocalMux t3727 (
    .I(seg_21_17_lutff_0_out_80932),
    .O(seg_21_17_local_g1_0_84812)
  );
  LocalMux t3728 (
    .I(seg_21_17_lutff_1_out_80933),
    .O(seg_21_17_local_g1_1_84813)
  );
  LocalMux t3729 (
    .I(seg_21_17_lutff_2_out_80934),
    .O(seg_21_17_local_g0_2_84806)
  );
  CascadeMux t373 (
    .I(net_56827),
    .O(net_56827_cascademuxed)
  );
  LocalMux t3730 (
    .I(seg_21_17_lutff_3_out_80935),
    .O(seg_21_17_local_g1_3_84815)
  );
  LocalMux t3731 (
    .I(seg_22_17_neigh_op_lft_3_80935),
    .O(seg_22_17_local_g0_3_88638)
  );
  LocalMux t3732 (
    .I(seg_20_17_neigh_op_rgt_4_80936),
    .O(seg_20_17_local_g3_4_81001)
  );
  LocalMux t3733 (
    .I(seg_22_17_neigh_op_lft_4_80936),
    .O(seg_22_17_local_g0_4_88639)
  );
  LocalMux t3734 (
    .I(seg_21_16_neigh_op_top_5_80937),
    .O(seg_21_16_local_g0_5_84686)
  );
  LocalMux t3735 (
    .I(seg_21_17_lutff_5_out_80937),
    .O(seg_21_17_local_g1_5_84817)
  );
  LocalMux t3736 (
    .I(seg_22_17_neigh_op_lft_5_80937),
    .O(seg_22_17_local_g0_5_88640)
  );
  LocalMux t3737 (
    .I(seg_20_17_neigh_op_rgt_6_80938),
    .O(seg_20_17_local_g3_6_81003)
  );
  LocalMux t3738 (
    .I(seg_20_18_neigh_op_bnr_6_80938),
    .O(seg_20_18_local_g0_6_81102)
  );
  LocalMux t3739 (
    .I(seg_22_16_neigh_op_tnl_6_80938),
    .O(seg_22_16_local_g2_6_88534)
  );
  CascadeMux t374 (
    .I(net_56839),
    .O(net_56839_cascademuxed)
  );
  LocalMux t3740 (
    .I(seg_21_17_lutff_7_out_80939),
    .O(seg_21_17_local_g3_7_84835)
  );
  LocalMux t3741 (
    .I(seg_22_17_neigh_op_lft_7_80939),
    .O(seg_22_17_local_g0_7_88642)
  );
  LocalMux t3742 (
    .I(seg_20_15_sp4_v_b_25_77215),
    .O(seg_20_15_local_g2_1_80744)
  );
  Span4Mux_v4 t3743 (
    .I(seg_20_17_sp4_h_r_1_81068),
    .O(seg_20_15_sp4_v_b_25_77215)
  );
  LocalMux t3744 (
    .I(seg_20_15_sp4_v_b_25_77215),
    .O(seg_20_15_local_g3_1_80752)
  );
  LocalMux t3745 (
    .I(seg_17_15_sp4_r_v_b_26_69851),
    .O(seg_17_15_local_g1_2_69875)
  );
  Span4Mux_v4 t3746 (
    .I(seg_18_17_sp4_h_r_9_74047),
    .O(seg_17_15_sp4_r_v_b_26_69851)
  );
  LocalMux t3747 (
    .I(seg_17_17_sp4_r_v_b_9_69856),
    .O(seg_17_17_local_g2_1_70128)
  );
  Span4Mux_v4 t3748 (
    .I(seg_18_17_sp4_h_r_9_74047),
    .O(seg_17_17_sp4_r_v_b_9_69856)
  );
  LocalMux t3749 (
    .I(seg_18_14_sp4_v_b_39_69851),
    .O(seg_18_14_local_g3_7_73604)
  );
  CascadeMux t375 (
    .I(net_56845),
    .O(net_56845_cascademuxed)
  );
  Span4Mux_v4 t3750 (
    .I(seg_18_17_sp4_h_r_9_74047),
    .O(seg_18_14_sp4_v_b_39_69851)
  );
  LocalMux t3751 (
    .I(seg_22_14_sp4_h_r_5_88367),
    .O(seg_22_14_local_g1_5_88279)
  );
  Span4Mux_h4 t3752 (
    .I(seg_22_14_sp4_v_t_37_84665),
    .O(seg_22_14_sp4_h_r_5_88367)
  );
  LocalMux t3753 (
    .I(seg_17_13_sp4_v_b_18_65654),
    .O(seg_17_13_local_g1_2_69629)
  );
  Span4Mux_v4 t3754 (
    .I(seg_17_14_sp4_h_r_7_69845),
    .O(seg_17_13_sp4_v_b_18_65654)
  );
  Span4Mux_h4 t3755 (
    .I(seg_21_14_sp4_v_t_36_80833),
    .O(seg_17_14_sp4_h_r_7_69845)
  );
  LocalMux t3756 (
    .I(seg_18_14_sp4_h_r_18_69845),
    .O(seg_18_14_local_g0_2_73575)
  );
  Span4Mux_h4 t3757 (
    .I(seg_21_14_sp4_v_t_36_80833),
    .O(seg_18_14_sp4_h_r_18_69845)
  );
  LocalMux t3758 (
    .I(seg_18_18_sp4_h_r_19_70336),
    .O(seg_18_18_local_g1_3_74076)
  );
  Span4Mux_h4 t3759 (
    .I(seg_21_18_sp4_v_b_1_80833),
    .O(seg_18_18_sp4_h_r_19_70336)
  );
  CascadeMux t376 (
    .I(net_56932),
    .O(net_56932_cascademuxed)
  );
  LocalMux t3760 (
    .I(seg_20_12_sp4_r_v_b_25_80341),
    .O(seg_20_12_local_g0_1_80359)
  );
  Span4Mux_v4 t3761 (
    .I(seg_21_14_sp4_v_t_36_80833),
    .O(seg_20_12_sp4_r_v_b_25_80341)
  );
  LocalMux t3762 (
    .I(seg_20_13_sp4_r_v_b_12_80341),
    .O(seg_20_13_local_g2_4_80501)
  );
  Span4Mux_v4 t3763 (
    .I(seg_21_14_sp4_v_t_36_80833),
    .O(seg_20_13_sp4_r_v_b_12_80341)
  );
  LocalMux t3764 (
    .I(seg_21_13_sp4_v_b_12_80341),
    .O(seg_21_13_local_g0_4_84316)
  );
  Span4Mux_v4 t3765 (
    .I(seg_21_14_sp4_v_t_36_80833),
    .O(seg_21_13_sp4_v_b_12_80341)
  );
  LocalMux t3766 (
    .I(seg_21_18_lutff_1_out_81056),
    .O(seg_21_18_local_g1_1_84936)
  );
  LocalMux t3767 (
    .I(seg_21_18_lutff_3_out_81058),
    .O(seg_21_18_local_g0_3_84930)
  );
  LocalMux t3768 (
    .I(seg_21_18_lutff_4_out_81059),
    .O(seg_21_18_local_g3_4_84955)
  );
  LocalMux t3769 (
    .I(seg_21_18_lutff_6_out_81061),
    .O(seg_21_18_local_g3_6_84957)
  );
  CascadeMux t377 (
    .I(net_56938),
    .O(net_56938_cascademuxed)
  );
  LocalMux t3770 (
    .I(seg_18_18_sp12_h_r_3_70324),
    .O(seg_18_18_local_g0_3_74068)
  );
  LocalMux t3771 (
    .I(seg_21_14_sp4_h_r_3_84534),
    .O(seg_21_14_local_g1_3_84446)
  );
  Span4Mux_h4 t3772 (
    .I(seg_21_14_sp4_v_t_47_80844),
    .O(seg_21_14_sp4_h_r_3_84534)
  );
  LocalMux t3773 (
    .I(seg_21_14_sp4_v_b_14_80466),
    .O(seg_21_14_local_g0_6_84441)
  );
  Span4Mux_v4 t3774 (
    .I(seg_21_15_sp4_v_t_38_80958),
    .O(seg_21_14_sp4_v_b_14_80466)
  );
  LocalMux t3775 (
    .I(seg_21_15_sp4_v_b_41_80838),
    .O(seg_21_15_local_g2_1_84575)
  );
  LocalMux t3776 (
    .I(seg_21_18_neigh_op_top_2_81180),
    .O(seg_21_18_local_g0_2_84929)
  );
  LocalMux t3777 (
    .I(seg_20_17_sp4_r_v_b_30_80963),
    .O(seg_20_17_local_g1_6_80987)
  );
  LocalMux t3778 (
    .I(seg_22_9_lutff_1_out_83780),
    .O(seg_22_9_local_g0_1_87652)
  );
  LocalMux t3779 (
    .I(seg_23_9_neigh_op_lft_1_83780),
    .O(seg_23_9_local_g1_1_91491)
  );
  CascadeMux t378 (
    .I(net_56950),
    .O(net_56950_cascademuxed)
  );
  LocalMux t3780 (
    .I(seg_21_13_neigh_op_rgt_2_84273),
    .O(seg_21_13_local_g3_2_84338)
  );
  LocalMux t3781 (
    .I(seg_21_13_sp4_h_r_31_77110),
    .O(seg_21_13_local_g3_7_84343)
  );
  LocalMux t3782 (
    .I(seg_18_14_sp4_r_v_b_8_73319),
    .O(seg_18_14_local_g2_0_73589)
  );
  Span4Mux_v4 t3783 (
    .I(seg_19_14_sp4_h_r_3_77208),
    .O(seg_18_14_sp4_r_v_b_8_73319)
  );
  LocalMux t3784 (
    .I(seg_22_14_neigh_op_top_4_84521),
    .O(seg_22_14_local_g0_4_88270)
  );
  LocalMux t3785 (
    .I(seg_22_17_sp4_r_v_b_13_88496),
    .O(seg_22_17_local_g2_5_88656)
  );
  LocalMux t3786 (
    .I(seg_21_17_sp4_r_v_b_12_84664),
    .O(seg_21_17_local_g2_4_84824)
  );
  LocalMux t3787 (
    .I(seg_21_15_neigh_op_tnr_7_84647),
    .O(seg_21_15_local_g2_7_84581)
  );
  LocalMux t3788 (
    .I(seg_21_17_neigh_op_rgt_2_84765),
    .O(seg_21_17_local_g2_2_84822)
  );
  LocalMux t3789 (
    .I(seg_21_17_neigh_op_rgt_5_84768),
    .O(seg_21_17_local_g3_5_84833)
  );
  CascadeMux t379 (
    .I(net_56956),
    .O(net_56956_cascademuxed)
  );
  LocalMux t3790 (
    .I(seg_21_17_neigh_op_rgt_6_84769),
    .O(seg_21_17_local_g2_6_84826)
  );
  LocalMux t3791 (
    .I(seg_19_13_sp4_h_r_30_69721),
    .O(seg_19_13_local_g3_6_77057)
  );
  Span4Mux_h4 t3792 (
    .I(seg_21_13_sp4_v_t_43_80717),
    .O(seg_19_13_sp4_h_r_30_69721)
  );
  Span4Mux_v4 t3793 (
    .I(seg_21_17_sp4_h_r_1_84899),
    .O(seg_21_13_sp4_v_t_43_80717)
  );
  LocalMux t3794 (
    .I(seg_19_17_sp4_h_r_33_70216),
    .O(seg_19_17_local_g2_1_77452)
  );
  Span4Mux_h4 t3795 (
    .I(seg_21_17_sp4_h_r_1_84899),
    .O(seg_19_17_sp4_h_r_33_70216)
  );
  LocalMux t3796 (
    .I(seg_19_17_sp4_h_r_30_70213),
    .O(seg_19_17_local_g2_6_77457)
  );
  Span4Mux_h4 t3797 (
    .I(seg_21_17_sp4_h_r_3_84903),
    .O(seg_19_17_sp4_h_r_30_70213)
  );
  LocalMux t3798 (
    .I(seg_18_17_sp4_h_r_14_70210),
    .O(seg_18_17_local_g0_6_73948)
  );
  Span4Mux_h4 t3799 (
    .I(seg_21_17_sp4_h_r_7_84907),
    .O(seg_18_17_sp4_h_r_14_70210)
  );
  CascadeMux t38 (
    .I(net_21135),
    .O(net_21135_cascademuxed)
  );
  CascadeMux t380 (
    .I(net_56962),
    .O(net_56962_cascademuxed)
  );
  LocalMux t3800 (
    .I(seg_18_17_sp4_h_r_22_70208),
    .O(seg_18_17_local_g1_6_73956)
  );
  Span4Mux_h4 t3801 (
    .I(seg_21_17_sp4_h_r_11_84901),
    .O(seg_18_17_sp4_h_r_22_70208)
  );
  LocalMux t3802 (
    .I(seg_19_15_sp4_v_b_25_73679),
    .O(seg_19_15_local_g2_1_77248)
  );
  Span4Mux_v4 t3803 (
    .I(seg_19_17_sp4_h_r_1_77510),
    .O(seg_19_15_sp4_v_b_25_73679)
  );
  LocalMux t3804 (
    .I(seg_19_17_sp4_h_r_1_77510),
    .O(seg_19_17_local_g0_1_77436)
  );
  LocalMux t3805 (
    .I(seg_19_15_sp4_v_b_32_73688),
    .O(seg_19_15_local_g2_0_77247)
  );
  Span4Mux_v4 t3806 (
    .I(seg_19_17_sp4_h_r_3_77514),
    .O(seg_19_15_sp4_v_b_32_73688)
  );
  LocalMux t3807 (
    .I(seg_19_17_sp4_h_r_3_77514),
    .O(seg_19_17_local_g1_3_77446)
  );
  LocalMux t3808 (
    .I(seg_19_15_sp4_v_b_29_73683),
    .O(seg_19_15_local_g2_5_77252)
  );
  Span4Mux_v4 t3809 (
    .I(seg_19_17_sp4_h_r_5_77516),
    .O(seg_19_15_sp4_v_b_29_73683)
  );
  CascadeMux t381 (
    .I(net_56968),
    .O(net_56968_cascademuxed)
  );
  LocalMux t3810 (
    .I(seg_19_17_sp4_h_r_5_77516),
    .O(seg_19_17_local_g0_5_77440)
  );
  LocalMux t3811 (
    .I(seg_19_15_sp4_v_b_31_73685),
    .O(seg_19_15_local_g3_7_77262)
  );
  Span4Mux_v4 t3812 (
    .I(seg_19_17_sp4_h_r_7_77518),
    .O(seg_19_15_sp4_v_b_31_73685)
  );
  LocalMux t3813 (
    .I(seg_19_17_sp4_h_r_7_77518),
    .O(seg_19_17_local_g1_7_77450)
  );
  LocalMux t3814 (
    .I(seg_19_13_sp4_v_b_7_73193),
    .O(seg_19_13_local_g1_7_77042)
  );
  Span4Mux_v4 t3815 (
    .I(seg_19_13_sp4_v_t_41_73684),
    .O(seg_19_13_sp4_v_b_7_73193)
  );
  Span4Mux_v4 t3816 (
    .I(seg_19_17_sp4_h_r_11_77512),
    .O(seg_19_13_sp4_v_t_41_73684)
  );
  LocalMux t3817 (
    .I(seg_19_15_sp4_v_b_28_73684),
    .O(seg_19_15_local_g2_4_77251)
  );
  Span4Mux_v4 t3818 (
    .I(seg_19_17_sp4_h_r_11_77512),
    .O(seg_19_15_sp4_v_b_28_73684)
  );
  LocalMux t3819 (
    .I(seg_18_17_sp4_h_r_11_74039),
    .O(seg_18_17_local_g1_3_73953)
  );
  CascadeMux t382 (
    .I(net_57061),
    .O(net_57061_cascademuxed)
  );
  Span4Mux_h4 t3820 (
    .I(seg_22_17_sp4_h_r_8_88739),
    .O(seg_18_17_sp4_h_r_11_74039)
  );
  LocalMux t3821 (
    .I(seg_19_13_sp4_h_r_5_77108),
    .O(seg_19_13_local_g1_5_77040)
  );
  Span4Mux_h4 t3822 (
    .I(seg_23_13_sp4_v_t_46_88382),
    .O(seg_19_13_sp4_h_r_5_77108)
  );
  LocalMux t3823 (
    .I(seg_19_13_sp4_h_r_9_77112),
    .O(seg_19_13_local_g1_1_77036)
  );
  Span4Mux_h4 t3824 (
    .I(seg_23_13_sp4_v_t_38_88374),
    .O(seg_19_13_sp4_h_r_9_77112)
  );
  LocalMux t3825 (
    .I(seg_19_13_sp4_h_r_11_77104),
    .O(seg_19_13_local_g0_3_77030)
  );
  Span4Mux_h4 t3826 (
    .I(seg_23_13_sp4_v_t_40_88376),
    .O(seg_19_13_sp4_h_r_11_77104)
  );
  LocalMux t3827 (
    .I(seg_22_15_sp4_v_b_38_84666),
    .O(seg_22_15_local_g3_6_88419)
  );
  LocalMux t3828 (
    .I(seg_19_17_sp4_h_r_18_74045),
    .O(seg_19_17_local_g0_2_77437)
  );
  Span4Mux_h4 t3829 (
    .I(seg_22_17_sp4_v_b_2_84544),
    .O(seg_19_17_sp4_h_r_18_74045)
  );
  CascadeMux t383 (
    .I(net_57085),
    .O(net_57085_cascademuxed)
  );
  LocalMux t3830 (
    .I(seg_19_15_sp4_h_r_17_73796),
    .O(seg_19_15_local_g0_1_77232)
  );
  Span4Mux_h4 t3831 (
    .I(seg_22_15_sp4_v_t_41_84792),
    .O(seg_19_15_sp4_h_r_17_73796)
  );
  LocalMux t3832 (
    .I(seg_19_15_sp4_h_r_23_73792),
    .O(seg_19_15_local_g1_7_77246)
  );
  Span4Mux_h4 t3833 (
    .I(seg_22_15_sp4_v_t_47_84798),
    .O(seg_19_15_sp4_h_r_23_73792)
  );
  LocalMux t3834 (
    .I(seg_19_13_sp4_h_r_19_73552),
    .O(seg_19_13_local_g1_3_77038)
  );
  Span4Mux_h4 t3835 (
    .I(seg_22_13_sp4_v_t_43_84548),
    .O(seg_19_13_sp4_h_r_19_73552)
  );
  LocalMux t3836 (
    .I(seg_19_13_sp4_h_r_15_73548),
    .O(seg_19_13_local_g0_7_77034)
  );
  Span4Mux_h4 t3837 (
    .I(seg_22_13_sp4_v_t_45_84550),
    .O(seg_19_13_sp4_h_r_15_73548)
  );
  LocalMux t3838 (
    .I(seg_23_9_lutff_2_out_87612),
    .O(seg_23_9_local_g0_2_91484)
  );
  LocalMux t3839 (
    .I(seg_20_6_sp4_h_r_20_76398),
    .O(seg_20_6_local_g0_4_79624)
  );
  CascadeMux t384 (
    .I(net_57097),
    .O(net_57097_cascademuxed)
  );
  Span4Mux_h4 t3840 (
    .I(seg_23_6_sp4_v_t_38_87513),
    .O(seg_20_6_sp4_h_r_20_76398)
  );
  CascadeMux t385 (
    .I(net_57430),
    .O(net_57430_cascademuxed)
  );
  CascadeMux t386 (
    .I(net_57460),
    .O(net_57460_cascademuxed)
  );
  CascadeMux t387 (
    .I(net_57466),
    .O(net_57466_cascademuxed)
  );
  CascadeMux t388 (
    .I(net_57571),
    .O(net_57571_cascademuxed)
  );
  CascadeMux t389 (
    .I(net_57583),
    .O(net_57583_cascademuxed)
  );
  CascadeMux t39 (
    .I(net_21141),
    .O(net_21141_cascademuxed)
  );
  CascadeMux t390 (
    .I(net_57589),
    .O(net_57589_cascademuxed)
  );
  CascadeMux t391 (
    .I(net_57676),
    .O(net_57676_cascademuxed)
  );
  CascadeMux t392 (
    .I(net_57682),
    .O(net_57682_cascademuxed)
  );
  CascadeMux t393 (
    .I(net_57688),
    .O(net_57688_cascademuxed)
  );
  CascadeMux t394 (
    .I(net_57694),
    .O(net_57694_cascademuxed)
  );
  CascadeMux t395 (
    .I(net_57700),
    .O(net_57700_cascademuxed)
  );
  CascadeMux t396 (
    .I(net_57706),
    .O(net_57706_cascademuxed)
  );
  CascadeMux t397 (
    .I(net_57712),
    .O(net_57712_cascademuxed)
  );
  CascadeMux t398 (
    .I(net_57835),
    .O(net_57835_cascademuxed)
  );
  CascadeMux t4 (
    .I(net_12225),
    .O(net_12225_cascademuxed)
  );
  CascadeMux t40 (
    .I(net_21228),
    .O(net_21228_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t400 (
    .carryinitin(),
    .carryinitout(t399)
  );
  CascadeMux t401 (
    .I(net_57928),
    .O(net_57928_cascademuxed)
  );
  CascadeMux t402 (
    .I(net_57940),
    .O(net_57940_cascademuxed)
  );
  CascadeMux t403 (
    .I(net_57952),
    .O(net_57952_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b10)
  ) t404 (
    .carryinitin(net_61785),
    .carryinitout(net_61829)
  );
  CascadeMux t405 (
    .I(net_58039),
    .O(net_58039_cascademuxed)
  );
  CascadeMux t406 (
    .I(net_58051),
    .O(net_58051_cascademuxed)
  );
  CascadeMux t407 (
    .I(net_58057),
    .O(net_58057_cascademuxed)
  );
  CascadeMux t408 (
    .I(net_58081),
    .O(net_58081_cascademuxed)
  );
  CascadeMux t409 (
    .I(net_58168),
    .O(net_58168_cascademuxed)
  );
  CascadeMux t41 (
    .I(net_21234),
    .O(net_21234_cascademuxed)
  );
  CascadeMux t410 (
    .I(net_58174),
    .O(net_58174_cascademuxed)
  );
  CascadeMux t411 (
    .I(net_58180),
    .O(net_58180_cascademuxed)
  );
  CascadeMux t412 (
    .I(net_58186),
    .O(net_58186_cascademuxed)
  );
  CascadeMux t413 (
    .I(net_58192),
    .O(net_58192_cascademuxed)
  );
  CascadeMux t414 (
    .I(net_58198),
    .O(net_58198_cascademuxed)
  );
  CascadeMux t415 (
    .I(net_58285),
    .O(net_58285_cascademuxed)
  );
  CascadeMux t416 (
    .I(net_58291),
    .O(net_58291_cascademuxed)
  );
  CascadeMux t417 (
    .I(net_58297),
    .O(net_58297_cascademuxed)
  );
  CascadeMux t418 (
    .I(net_58309),
    .O(net_58309_cascademuxed)
  );
  CascadeMux t419 (
    .I(net_58315),
    .O(net_58315_cascademuxed)
  );
  CascadeMux t42 (
    .I(net_21246),
    .O(net_21246_cascademuxed)
  );
  CascadeMux t420 (
    .I(net_58327),
    .O(net_58327_cascademuxed)
  );
  CascadeMux t421 (
    .I(net_58414),
    .O(net_58414_cascademuxed)
  );
  CascadeMux t422 (
    .I(net_58420),
    .O(net_58420_cascademuxed)
  );
  CascadeMux t423 (
    .I(net_58426),
    .O(net_58426_cascademuxed)
  );
  CascadeMux t424 (
    .I(net_58432),
    .O(net_58432_cascademuxed)
  );
  CascadeMux t425 (
    .I(net_58438),
    .O(net_58438_cascademuxed)
  );
  CascadeMux t426 (
    .I(net_58531),
    .O(net_58531_cascademuxed)
  );
  CascadeMux t427 (
    .I(net_58537),
    .O(net_58537_cascademuxed)
  );
  CascadeMux t428 (
    .I(net_58555),
    .O(net_58555_cascademuxed)
  );
  CascadeMux t429 (
    .I(net_58801),
    .O(net_58801_cascademuxed)
  );
  CascadeMux t43 (
    .I(net_21351),
    .O(net_21351_cascademuxed)
  );
  CascadeMux t430 (
    .I(net_58819),
    .O(net_58819_cascademuxed)
  );
  CascadeMux t431 (
    .I(net_58906),
    .O(net_58906_cascademuxed)
  );
  CascadeMux t432 (
    .I(net_58936),
    .O(net_58936_cascademuxed)
  );
  CascadeMux t433 (
    .I(net_59023),
    .O(net_59023_cascademuxed)
  );
  CascadeMux t434 (
    .I(net_59029),
    .O(net_59029_cascademuxed)
  );
  CascadeMux t435 (
    .I(net_59035),
    .O(net_59035_cascademuxed)
  );
  CascadeMux t436 (
    .I(net_59053),
    .O(net_59053_cascademuxed)
  );
  CascadeMux t437 (
    .I(net_59065),
    .O(net_59065_cascademuxed)
  );
  CascadeMux t438 (
    .I(net_59785),
    .O(net_59785_cascademuxed)
  );
  CascadeMux t439 (
    .I(net_59890),
    .O(net_59890_cascademuxed)
  );
  CascadeMux t44 (
    .I(net_23331),
    .O(net_23331_cascademuxed)
  );
  CascadeMux t440 (
    .I(net_59914),
    .O(net_59914_cascademuxed)
  );
  CascadeMux t441 (
    .I(net_60639),
    .O(net_60639_cascademuxed)
  );
  CascadeMux t442 (
    .I(net_60645),
    .O(net_60645_cascademuxed)
  );
  CascadeMux t443 (
    .I(net_60651),
    .O(net_60651_cascademuxed)
  );
  CascadeMux t444 (
    .I(net_60657),
    .O(net_60657_cascademuxed)
  );
  CascadeMux t445 (
    .I(net_60768),
    .O(net_60768_cascademuxed)
  );
  CascadeMux t446 (
    .I(net_60786),
    .O(net_60786_cascademuxed)
  );
  CascadeMux t447 (
    .I(net_60792),
    .O(net_60792_cascademuxed)
  );
  CascadeMux t448 (
    .I(net_60798),
    .O(net_60798_cascademuxed)
  );
  CascadeMux t449 (
    .I(net_60804),
    .O(net_60804_cascademuxed)
  );
  CascadeMux t45 (
    .I(net_25188),
    .O(net_25188_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t451 (
    .carryinitin(),
    .carryinitout(t450)
  );
  CascadeMux t453 (
    .I(net_61530),
    .O(net_61530_cascademuxed)
  );
  CascadeMux t454 (
    .I(net_61542),
    .O(net_61542_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t456 (
    .carryinitin(),
    .carryinitout(t455)
  );
  CascadeMux t457 (
    .I(net_61623),
    .O(net_61623_cascademuxed)
  );
  CascadeMux t459 (
    .I(net_61629),
    .O(net_61629_cascademuxed)
  );
  CascadeMux t460 (
    .I(net_61647),
    .O(net_61647_cascademuxed)
  );
  CascadeMux t461 (
    .I(net_61653),
    .O(net_61653_cascademuxed)
  );
  CascadeMux t462 (
    .I(net_61659),
    .O(net_61659_cascademuxed)
  );
  CascadeMux t463 (
    .I(net_61746),
    .O(net_61746_cascademuxed)
  );
  CascadeMux t464 (
    .I(net_61752),
    .O(net_61752_cascademuxed)
  );
  CascadeMux t465 (
    .I(net_61758),
    .O(net_61758_cascademuxed)
  );
  CascadeMux t466 (
    .I(net_61764),
    .O(net_61764_cascademuxed)
  );
  CascadeMux t467 (
    .I(net_61770),
    .O(net_61770_cascademuxed)
  );
  CascadeMux t468 (
    .I(net_61776),
    .O(net_61776_cascademuxed)
  );
  CascadeMux t469 (
    .I(net_61782),
    .O(net_61782_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t47 (
    .carryinitin(),
    .carryinitout(t46)
  );
  CascadeMux t470 (
    .I(net_61788),
    .O(net_61788_cascademuxed)
  );
  CascadeMux t471 (
    .I(net_61869),
    .O(net_61869_cascademuxed)
  );
  CascadeMux t472 (
    .I(net_61875),
    .O(net_61875_cascademuxed)
  );
  CascadeMux t473 (
    .I(net_61881),
    .O(net_61881_cascademuxed)
  );
  CascadeMux t474 (
    .I(net_61887),
    .O(net_61887_cascademuxed)
  );
  CascadeMux t475 (
    .I(net_61893),
    .O(net_61893_cascademuxed)
  );
  CascadeMux t476 (
    .I(net_61899),
    .O(net_61899_cascademuxed)
  );
  CascadeMux t477 (
    .I(net_61905),
    .O(net_61905_cascademuxed)
  );
  CascadeMux t478 (
    .I(net_61911),
    .O(net_61911_cascademuxed)
  );
  CascadeMux t479 (
    .I(net_61992),
    .O(net_61992_cascademuxed)
  );
  CascadeMux t480 (
    .I(net_61998),
    .O(net_61998_cascademuxed)
  );
  CascadeMux t481 (
    .I(net_62004),
    .O(net_62004_cascademuxed)
  );
  CascadeMux t482 (
    .I(net_62010),
    .O(net_62010_cascademuxed)
  );
  CascadeMux t483 (
    .I(net_62022),
    .O(net_62022_cascademuxed)
  );
  CascadeMux t484 (
    .I(net_62028),
    .O(net_62028_cascademuxed)
  );
  CascadeMux t485 (
    .I(net_62034),
    .O(net_62034_cascademuxed)
  );
  CascadeMux t486 (
    .I(net_62121),
    .O(net_62121_cascademuxed)
  );
  CascadeMux t487 (
    .I(net_62139),
    .O(net_62139_cascademuxed)
  );
  CascadeMux t488 (
    .I(net_62145),
    .O(net_62145_cascademuxed)
  );
  CascadeMux t489 (
    .I(net_62157),
    .O(net_62157_cascademuxed)
  );
  CascadeMux t49 (
    .I(net_29836),
    .O(net_29836_cascademuxed)
  );
  CascadeMux t490 (
    .I(net_62250),
    .O(net_62250_cascademuxed)
  );
  CascadeMux t491 (
    .I(net_62256),
    .O(net_62256_cascademuxed)
  );
  CascadeMux t492 (
    .I(net_62262),
    .O(net_62262_cascademuxed)
  );
  CascadeMux t493 (
    .I(net_62268),
    .O(net_62268_cascademuxed)
  );
  CascadeMux t494 (
    .I(net_62280),
    .O(net_62280_cascademuxed)
  );
  CascadeMux t495 (
    .I(net_62385),
    .O(net_62385_cascademuxed)
  );
  CascadeMux t496 (
    .I(net_62403),
    .O(net_62403_cascademuxed)
  );
  CascadeMux t497 (
    .I(net_62484),
    .O(net_62484_cascademuxed)
  );
  CascadeMux t498 (
    .I(net_62490),
    .O(net_62490_cascademuxed)
  );
  CascadeMux t499 (
    .I(net_62502),
    .O(net_62502_cascademuxed)
  );
  CascadeMux t5 (
    .I(net_12231),
    .O(net_12231_cascademuxed)
  );
  CascadeMux t500 (
    .I(net_62526),
    .O(net_62526_cascademuxed)
  );
  CascadeMux t501 (
    .I(net_62607),
    .O(net_62607_cascademuxed)
  );
  CascadeMux t502 (
    .I(net_62613),
    .O(net_62613_cascademuxed)
  );
  CascadeMux t503 (
    .I(net_62619),
    .O(net_62619_cascademuxed)
  );
  CascadeMux t504 (
    .I(net_62643),
    .O(net_62643_cascademuxed)
  );
  CascadeMux t505 (
    .I(net_62748),
    .O(net_62748_cascademuxed)
  );
  CascadeMux t506 (
    .I(net_62766),
    .O(net_62766_cascademuxed)
  );
  CascadeMux t507 (
    .I(net_62865),
    .O(net_62865_cascademuxed)
  );
  CascadeMux t508 (
    .I(net_62889),
    .O(net_62889_cascademuxed)
  );
  CascadeMux t509 (
    .I(net_62895),
    .O(net_62895_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t51 (
    .carryinitin(),
    .carryinitout(t50)
  );
  CascadeMux t510 (
    .I(net_63228),
    .O(net_63228_cascademuxed)
  );
  CascadeMux t511 (
    .I(net_63252),
    .O(net_63252_cascademuxed)
  );
  CascadeMux t512 (
    .I(net_63264),
    .O(net_63264_cascademuxed)
  );
  CascadeMux t513 (
    .I(net_63837),
    .O(net_63837_cascademuxed)
  );
  CascadeMux t514 (
    .I(net_63861),
    .O(net_63861_cascademuxed)
  );
  CascadeMux t515 (
    .I(net_63867),
    .O(net_63867_cascademuxed)
  );
  CascadeMux t516 (
    .I(net_63879),
    .O(net_63879_cascademuxed)
  );
  CascadeMux t517 (
    .I(net_63990),
    .O(net_63990_cascademuxed)
  );
  CascadeMux t518 (
    .I(net_64002),
    .O(net_64002_cascademuxed)
  );
  CascadeMux t519 (
    .I(net_64488),
    .O(net_64488_cascademuxed)
  );
  CascadeMux t520 (
    .I(net_64500),
    .O(net_64500_cascademuxed)
  );
  CascadeMux t521 (
    .I(net_64845),
    .O(net_64845_cascademuxed)
  );
  CascadeMux t522 (
    .I(net_64962),
    .O(net_64962_cascademuxed)
  );
  CascadeMux t523 (
    .I(net_65343),
    .O(net_65343_cascademuxed)
  );
  CascadeMux t524 (
    .I(net_65355),
    .O(net_65355_cascademuxed)
  );
  CascadeMux t525 (
    .I(net_65361),
    .O(net_65361_cascademuxed)
  );
  CascadeMux t526 (
    .I(net_65367),
    .O(net_65367_cascademuxed)
  );
  CascadeMux t527 (
    .I(net_65583),
    .O(net_65583_cascademuxed)
  );
  CascadeMux t528 (
    .I(net_65700),
    .O(net_65700_cascademuxed)
  );
  CascadeMux t529 (
    .I(net_65706),
    .O(net_65706_cascademuxed)
  );
  CascadeMux t53 (
    .I(net_31223),
    .O(net_31223_cascademuxed)
  );
  CascadeMux t530 (
    .I(net_65712),
    .O(net_65712_cascademuxed)
  );
  CascadeMux t531 (
    .I(net_65730),
    .O(net_65730_cascademuxed)
  );
  CascadeMux t532 (
    .I(net_65736),
    .O(net_65736_cascademuxed)
  );
  CascadeMux t533 (
    .I(net_65835),
    .O(net_65835_cascademuxed)
  );
  CascadeMux t534 (
    .I(net_65952),
    .O(net_65952_cascademuxed)
  );
  CascadeMux t535 (
    .I(net_65976),
    .O(net_65976_cascademuxed)
  );
  CascadeMux t536 (
    .I(net_66069),
    .O(net_66069_cascademuxed)
  );
  CascadeMux t537 (
    .I(net_66081),
    .O(net_66081_cascademuxed)
  );
  CascadeMux t538 (
    .I(net_66087),
    .O(net_66087_cascademuxed)
  );
  CascadeMux t539 (
    .I(net_66099),
    .O(net_66099_cascademuxed)
  );
  CascadeMux t54 (
    .I(net_31253),
    .O(net_31253_cascademuxed)
  );
  CascadeMux t540 (
    .I(net_66105),
    .O(net_66105_cascademuxed)
  );
  CascadeMux t541 (
    .I(net_66198),
    .O(net_66198_cascademuxed)
  );
  CascadeMux t542 (
    .I(net_66321),
    .O(net_66321_cascademuxed)
  );
  CascadeMux t543 (
    .I(net_66450),
    .O(net_66450_cascademuxed)
  );
  CascadeMux t544 (
    .I(net_66456),
    .O(net_66456_cascademuxed)
  );
  CascadeMux t545 (
    .I(net_66567),
    .O(net_66567_cascademuxed)
  );
  CascadeMux t546 (
    .I(net_66585),
    .O(net_66585_cascademuxed)
  );
  CascadeMux t547 (
    .I(net_66591),
    .O(net_66591_cascademuxed)
  );
  CascadeMux t548 (
    .I(net_66597),
    .O(net_66597_cascademuxed)
  );
  CascadeMux t549 (
    .I(net_66690),
    .O(net_66690_cascademuxed)
  );
  CascadeMux t550 (
    .I(net_66696),
    .O(net_66696_cascademuxed)
  );
  CascadeMux t551 (
    .I(net_66702),
    .O(net_66702_cascademuxed)
  );
  CascadeMux t552 (
    .I(net_66708),
    .O(net_66708_cascademuxed)
  );
  CascadeMux t553 (
    .I(net_66714),
    .O(net_66714_cascademuxed)
  );
  CascadeMux t554 (
    .I(net_67674),
    .O(net_67674_cascademuxed)
  );
  CascadeMux t555 (
    .I(net_67680),
    .O(net_67680_cascademuxed)
  );
  CascadeMux t556 (
    .I(net_67686),
    .O(net_67686_cascademuxed)
  );
  CascadeMux t557 (
    .I(net_67698),
    .O(net_67698_cascademuxed)
  );
  CascadeMux t558 (
    .I(net_67704),
    .O(net_67704_cascademuxed)
  );
  CascadeMux t559 (
    .I(net_67710),
    .O(net_67710_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t56 (
    .carryinitin(),
    .carryinitout(t55)
  );
  CascadeMux t560 (
    .I(net_67791),
    .O(net_67791_cascademuxed)
  );
  CascadeMux t561 (
    .I(net_67815),
    .O(net_67815_cascademuxed)
  );
  CascadeMux t562 (
    .I(net_67827),
    .O(net_67827_cascademuxed)
  );
  CascadeMux t563 (
    .I(net_68670),
    .O(net_68670_cascademuxed)
  );
  CascadeMux t564 (
    .I(net_68706),
    .O(net_68706_cascademuxed)
  );
  CascadeMux t565 (
    .I(net_68712),
    .O(net_68712_cascademuxed)
  );
  CascadeMux t566 (
    .I(net_68817),
    .O(net_68817_cascademuxed)
  );
  CascadeMux t567 (
    .I(net_68823),
    .O(net_68823_cascademuxed)
  );
  CascadeMux t568 (
    .I(net_68835),
    .O(net_68835_cascademuxed)
  );
  CascadeMux t569 (
    .I(net_69690),
    .O(net_69690_cascademuxed)
  );
  CascadeMux t570 (
    .I(net_69807),
    .O(net_69807_cascademuxed)
  );
  CascadeMux t571 (
    .I(net_69900),
    .O(net_69900_cascademuxed)
  );
  CascadeMux t572 (
    .I(net_69918),
    .O(net_69918_cascademuxed)
  );
  CascadeMux t573 (
    .I(net_69924),
    .O(net_69924_cascademuxed)
  );
  CascadeMux t574 (
    .I(net_70065),
    .O(net_70065_cascademuxed)
  );
  CascadeMux t575 (
    .I(net_70146),
    .O(net_70146_cascademuxed)
  );
  CascadeMux t576 (
    .I(net_70158),
    .O(net_70158_cascademuxed)
  );
  CascadeMux t577 (
    .I(net_70176),
    .O(net_70176_cascademuxed)
  );
  CascadeMux t578 (
    .I(net_70188),
    .O(net_70188_cascademuxed)
  );
  CascadeMux t579 (
    .I(net_70269),
    .O(net_70269_cascademuxed)
  );
  CascadeMux t58 (
    .I(net_33830),
    .O(net_33830_cascademuxed)
  );
  CascadeMux t580 (
    .I(net_70293),
    .O(net_70293_cascademuxed)
  );
  CascadeMux t581 (
    .I(net_70305),
    .O(net_70305_cascademuxed)
  );
  CascadeMux t582 (
    .I(net_70398),
    .O(net_70398_cascademuxed)
  );
  CascadeMux t583 (
    .I(net_70416),
    .O(net_70416_cascademuxed)
  );
  CascadeMux t584 (
    .I(net_70428),
    .O(net_70428_cascademuxed)
  );
  CascadeMux t585 (
    .I(net_70434),
    .O(net_70434_cascademuxed)
  );
  CascadeMux t586 (
    .I(net_70515),
    .O(net_70515_cascademuxed)
  );
  CascadeMux t587 (
    .I(net_70521),
    .O(net_70521_cascademuxed)
  );
  CascadeMux t588 (
    .I(net_70668),
    .O(net_70668_cascademuxed)
  );
  CascadeMux t589 (
    .I(net_71652),
    .O(net_71652_cascademuxed)
  );
  CascadeMux t59 (
    .I(net_33842),
    .O(net_33842_cascademuxed)
  );
  CascadeMux t590 (
    .I(net_71658),
    .O(net_71658_cascademuxed)
  );
  CascadeMux t591 (
    .I(net_71664),
    .O(net_71664_cascademuxed)
  );
  CascadeMux t592 (
    .I(net_72624),
    .O(net_72624_cascademuxed)
  );
  CascadeMux t593 (
    .I(net_72630),
    .O(net_72630_cascademuxed)
  );
  CascadeMux t594 (
    .I(net_72654),
    .O(net_72654_cascademuxed)
  );
  CascadeMux t595 (
    .I(net_72660),
    .O(net_72660_cascademuxed)
  );
  CascadeMux t596 (
    .I(net_72666),
    .O(net_72666_cascademuxed)
  );
  CascadeMux t597 (
    .I(net_73134),
    .O(net_73134_cascademuxed)
  );
  CascadeMux t598 (
    .I(net_73497),
    .O(net_73497_cascademuxed)
  );
  CascadeMux t599 (
    .I(net_73503),
    .O(net_73503_cascademuxed)
  );
  CascadeMux t6 (
    .I(net_12243),
    .O(net_12243_cascademuxed)
  );
  CascadeMux t60 (
    .I(net_33848),
    .O(net_33848_cascademuxed)
  );
  CascadeMux t600 (
    .I(net_73509),
    .O(net_73509_cascademuxed)
  );
  CascadeMux t601 (
    .I(net_73527),
    .O(net_73527_cascademuxed)
  );
  CascadeMux t602 (
    .I(net_73608),
    .O(net_73608_cascademuxed)
  );
  CascadeMux t603 (
    .I(net_73614),
    .O(net_73614_cascademuxed)
  );
  CascadeMux t604 (
    .I(net_73632),
    .O(net_73632_cascademuxed)
  );
  CascadeMux t605 (
    .I(net_73650),
    .O(net_73650_cascademuxed)
  );
  CascadeMux t606 (
    .I(net_73749),
    .O(net_73749_cascademuxed)
  );
  CascadeMux t607 (
    .I(net_73767),
    .O(net_73767_cascademuxed)
  );
  CascadeMux t608 (
    .I(net_73983),
    .O(net_73983_cascademuxed)
  );
  CascadeMux t609 (
    .I(net_74001),
    .O(net_74001_cascademuxed)
  );
  CascadeMux t61 (
    .I(net_33854),
    .O(net_33854_cascademuxed)
  );
  CascadeMux t610 (
    .I(net_74007),
    .O(net_74007_cascademuxed)
  );
  CascadeMux t611 (
    .I(net_74013),
    .O(net_74013_cascademuxed)
  );
  CascadeMux t612 (
    .I(net_74112),
    .O(net_74112_cascademuxed)
  );
  CascadeMux t613 (
    .I(net_74124),
    .O(net_74124_cascademuxed)
  );
  CascadeMux t614 (
    .I(net_77075),
    .O(net_77075_cascademuxed)
  );
  CascadeMux t615 (
    .I(net_77076),
    .O(net_77076_cascademuxed)
  );
  CascadeMux t616 (
    .I(net_77078),
    .O(net_77078_cascademuxed)
  );
  CascadeMux t617 (
    .I(net_77079),
    .O(net_77079_cascademuxed)
  );
  CascadeMux t618 (
    .I(net_77080),
    .O(net_77080_cascademuxed)
  );
  CascadeMux t619 (
    .I(net_77081),
    .O(net_77081_cascademuxed)
  );
  CascadeMux t62 (
    .I(net_33860),
    .O(net_33860_cascademuxed)
  );
  CascadeMux t620 (
    .I(net_77082),
    .O(net_77082_cascademuxed)
  );
  CascadeMux t621 (
    .I(net_77083),
    .O(net_77083_cascademuxed)
  );
  CascadeMux t622 (
    .I(net_77177),
    .O(net_77177_cascademuxed)
  );
  CascadeMux t623 (
    .I(net_77178),
    .O(net_77178_cascademuxed)
  );
  CascadeMux t624 (
    .I(net_77180),
    .O(net_77180_cascademuxed)
  );
  CascadeMux t625 (
    .I(net_77181),
    .O(net_77181_cascademuxed)
  );
  CascadeMux t626 (
    .I(net_77182),
    .O(net_77182_cascademuxed)
  );
  CascadeMux t627 (
    .I(net_77183),
    .O(net_77183_cascademuxed)
  );
  CascadeMux t628 (
    .I(net_77184),
    .O(net_77184_cascademuxed)
  );
  CascadeMux t629 (
    .I(net_77185),
    .O(net_77185_cascademuxed)
  );
  CascadeMux t63 (
    .I(net_33866),
    .O(net_33866_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t631 (
    .carryinitin(),
    .carryinitout(t630)
  );
  CascadeMux t632 (
    .I(net_77279),
    .O(net_77279_cascademuxed)
  );
  CascadeMux t633 (
    .I(net_77280),
    .O(net_77280_cascademuxed)
  );
  CascadeMux t634 (
    .I(net_77282),
    .O(net_77282_cascademuxed)
  );
  CascadeMux t635 (
    .I(net_77283),
    .O(net_77283_cascademuxed)
  );
  CascadeMux t636 (
    .I(net_77284),
    .O(net_77284_cascademuxed)
  );
  CascadeMux t637 (
    .I(net_77285),
    .O(net_77285_cascademuxed)
  );
  CascadeMux t638 (
    .I(net_77286),
    .O(net_77286_cascademuxed)
  );
  CascadeMux t639 (
    .I(net_77287),
    .O(net_77287_cascademuxed)
  );
  CascadeMux t64 (
    .I(net_33971),
    .O(net_33971_cascademuxed)
  );
  CascadeMux t640 (
    .I(net_77381),
    .O(net_77381_cascademuxed)
  );
  CascadeMux t641 (
    .I(net_77382),
    .O(net_77382_cascademuxed)
  );
  CascadeMux t642 (
    .I(net_77384),
    .O(net_77384_cascademuxed)
  );
  CascadeMux t643 (
    .I(net_77385),
    .O(net_77385_cascademuxed)
  );
  CascadeMux t644 (
    .I(net_77386),
    .O(net_77386_cascademuxed)
  );
  CascadeMux t645 (
    .I(net_77387),
    .O(net_77387_cascademuxed)
  );
  CascadeMux t646 (
    .I(net_77388),
    .O(net_77388_cascademuxed)
  );
  CascadeMux t647 (
    .I(net_77389),
    .O(net_77389_cascademuxed)
  );
  CascadeMux t648 (
    .I(net_77483),
    .O(net_77483_cascademuxed)
  );
  CascadeMux t649 (
    .I(net_77484),
    .O(net_77484_cascademuxed)
  );
  CascadeMux t65 (
    .I(net_33977),
    .O(net_33977_cascademuxed)
  );
  CascadeMux t650 (
    .I(net_77486),
    .O(net_77486_cascademuxed)
  );
  CascadeMux t651 (
    .I(net_77487),
    .O(net_77487_cascademuxed)
  );
  CascadeMux t652 (
    .I(net_77488),
    .O(net_77488_cascademuxed)
  );
  CascadeMux t653 (
    .I(net_77489),
    .O(net_77489_cascademuxed)
  );
  CascadeMux t654 (
    .I(net_77490),
    .O(net_77490_cascademuxed)
  );
  CascadeMux t655 (
    .I(net_77491),
    .O(net_77491_cascademuxed)
  );
  CascadeMux t656 (
    .I(net_77585),
    .O(net_77585_cascademuxed)
  );
  CascadeMux t657 (
    .I(net_77586),
    .O(net_77586_cascademuxed)
  );
  CascadeMux t658 (
    .I(net_77588),
    .O(net_77588_cascademuxed)
  );
  CascadeMux t659 (
    .I(net_77589),
    .O(net_77589_cascademuxed)
  );
  CascadeMux t66 (
    .I(net_33983),
    .O(net_33983_cascademuxed)
  );
  CascadeMux t660 (
    .I(net_77590),
    .O(net_77590_cascademuxed)
  );
  CascadeMux t661 (
    .I(net_77591),
    .O(net_77591_cascademuxed)
  );
  CascadeMux t662 (
    .I(net_77592),
    .O(net_77592_cascademuxed)
  );
  CascadeMux t663 (
    .I(net_77593),
    .O(net_77593_cascademuxed)
  );
  CascadeMux t664 (
    .I(net_79655),
    .O(net_79655_cascademuxed)
  );
  CascadeMux t665 (
    .I(net_79667),
    .O(net_79667_cascademuxed)
  );
  CascadeMux t666 (
    .I(net_79685),
    .O(net_79685_cascademuxed)
  );
  CascadeMux t667 (
    .I(net_79697),
    .O(net_79697_cascademuxed)
  );
  CascadeMux t668 (
    .I(net_79778),
    .O(net_79778_cascademuxed)
  );
  CascadeMux t669 (
    .I(net_80147),
    .O(net_80147_cascademuxed)
  );
  CascadeMux t670 (
    .I(net_80165),
    .O(net_80165_cascademuxed)
  );
  CascadeMux t671 (
    .I(net_80177),
    .O(net_80177_cascademuxed)
  );
  CascadeMux t672 (
    .I(net_80189),
    .O(net_80189_cascademuxed)
  );
  CascadeMux t673 (
    .I(net_80300),
    .O(net_80300_cascademuxed)
  );
  CascadeMux t674 (
    .I(net_80393),
    .O(net_80393_cascademuxed)
  );
  CascadeMux t675 (
    .I(net_80405),
    .O(net_80405_cascademuxed)
  );
  CascadeMux t676 (
    .I(net_80417),
    .O(net_80417_cascademuxed)
  );
  CascadeMux t677 (
    .I(net_80429),
    .O(net_80429_cascademuxed)
  );
  CascadeMux t678 (
    .I(net_80435),
    .O(net_80435_cascademuxed)
  );
  CascadeMux t679 (
    .I(net_80516),
    .O(net_80516_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t68 (
    .carryinitin(),
    .carryinitout(t67)
  );
  CascadeMux t680 (
    .I(net_80522),
    .O(net_80522_cascademuxed)
  );
  CascadeMux t681 (
    .I(net_80528),
    .O(net_80528_cascademuxed)
  );
  CascadeMux t682 (
    .I(net_80540),
    .O(net_80540_cascademuxed)
  );
  CascadeMux t683 (
    .I(net_80552),
    .O(net_80552_cascademuxed)
  );
  CascadeMux t684 (
    .I(net_80558),
    .O(net_80558_cascademuxed)
  );
  CascadeMux t685 (
    .I(net_80639),
    .O(net_80639_cascademuxed)
  );
  CascadeMux t686 (
    .I(net_80657),
    .O(net_80657_cascademuxed)
  );
  CascadeMux t687 (
    .I(net_80669),
    .O(net_80669_cascademuxed)
  );
  CascadeMux t688 (
    .I(net_80681),
    .O(net_80681_cascademuxed)
  );
  CascadeMux t689 (
    .I(net_80762),
    .O(net_80762_cascademuxed)
  );
  CascadeMux t690 (
    .I(net_80768),
    .O(net_80768_cascademuxed)
  );
  CascadeMux t691 (
    .I(net_80774),
    .O(net_80774_cascademuxed)
  );
  CascadeMux t692 (
    .I(net_80780),
    .O(net_80780_cascademuxed)
  );
  CascadeMux t693 (
    .I(net_80798),
    .O(net_80798_cascademuxed)
  );
  CascadeMux t694 (
    .I(net_80804),
    .O(net_80804_cascademuxed)
  );
  CascadeMux t695 (
    .I(net_80885),
    .O(net_80885_cascademuxed)
  );
  CascadeMux t696 (
    .I(net_80897),
    .O(net_80897_cascademuxed)
  );
  CascadeMux t697 (
    .I(net_80915),
    .O(net_80915_cascademuxed)
  );
  CascadeMux t698 (
    .I(net_81008),
    .O(net_81008_cascademuxed)
  );
  CascadeMux t699 (
    .I(net_81014),
    .O(net_81014_cascademuxed)
  );
  CascadeMux t7 (
    .I(net_12249),
    .O(net_12249_cascademuxed)
  );
  CascadeMux t70 (
    .I(net_34820),
    .O(net_34820_cascademuxed)
  );
  CascadeMux t700 (
    .I(net_81020),
    .O(net_81020_cascademuxed)
  );
  CascadeMux t701 (
    .I(net_81032),
    .O(net_81032_cascademuxed)
  );
  CascadeMux t702 (
    .I(net_81038),
    .O(net_81038_cascademuxed)
  );
  CascadeMux t703 (
    .I(net_81044),
    .O(net_81044_cascademuxed)
  );
  CascadeMux t704 (
    .I(net_81050),
    .O(net_81050_cascademuxed)
  );
  CascadeMux t705 (
    .I(net_81149),
    .O(net_81149_cascademuxed)
  );
  CascadeMux t706 (
    .I(net_81155),
    .O(net_81155_cascademuxed)
  );
  CascadeMux t707 (
    .I(net_81161),
    .O(net_81161_cascademuxed)
  );
  CascadeMux t708 (
    .I(net_81173),
    .O(net_81173_cascademuxed)
  );
  CascadeMux t709 (
    .I(net_83504),
    .O(net_83504_cascademuxed)
  );
  CascadeMux t71 (
    .I(net_34838),
    .O(net_34838_cascademuxed)
  );
  CascadeMux t710 (
    .I(net_83855),
    .O(net_83855_cascademuxed)
  );
  CascadeMux t711 (
    .I(net_83867),
    .O(net_83867_cascademuxed)
  );
  CascadeMux t712 (
    .I(net_83978),
    .O(net_83978_cascademuxed)
  );
  CascadeMux t713 (
    .I(net_84002),
    .O(net_84002_cascademuxed)
  );
  CascadeMux t714 (
    .I(net_84254),
    .O(net_84254_cascademuxed)
  );
  CascadeMux t715 (
    .I(net_84347),
    .O(net_84347_cascademuxed)
  );
  CascadeMux t716 (
    .I(net_84353),
    .O(net_84353_cascademuxed)
  );
  CascadeMux t717 (
    .I(net_84359),
    .O(net_84359_cascademuxed)
  );
  CascadeMux t718 (
    .I(net_84371),
    .O(net_84371_cascademuxed)
  );
  CascadeMux t719 (
    .I(net_84383),
    .O(net_84383_cascademuxed)
  );
  CascadeMux t72 (
    .I(net_34844),
    .O(net_34844_cascademuxed)
  );
  CascadeMux t720 (
    .I(net_84476),
    .O(net_84476_cascademuxed)
  );
  CascadeMux t721 (
    .I(net_84482),
    .O(net_84482_cascademuxed)
  );
  CascadeMux t722 (
    .I(net_84488),
    .O(net_84488_cascademuxed)
  );
  CascadeMux t723 (
    .I(net_84494),
    .O(net_84494_cascademuxed)
  );
  CascadeMux t724 (
    .I(net_84500),
    .O(net_84500_cascademuxed)
  );
  CascadeMux t725 (
    .I(net_84506),
    .O(net_84506_cascademuxed)
  );
  CascadeMux t726 (
    .I(net_84512),
    .O(net_84512_cascademuxed)
  );
  CascadeMux t727 (
    .I(net_84593),
    .O(net_84593_cascademuxed)
  );
  CascadeMux t728 (
    .I(net_84599),
    .O(net_84599_cascademuxed)
  );
  CascadeMux t729 (
    .I(net_84605),
    .O(net_84605_cascademuxed)
  );
  CascadeMux t73 (
    .I(net_34850),
    .O(net_34850_cascademuxed)
  );
  CascadeMux t730 (
    .I(net_84617),
    .O(net_84617_cascademuxed)
  );
  CascadeMux t731 (
    .I(net_84623),
    .O(net_84623_cascademuxed)
  );
  CascadeMux t732 (
    .I(net_84629),
    .O(net_84629_cascademuxed)
  );
  CascadeMux t733 (
    .I(net_84635),
    .O(net_84635_cascademuxed)
  );
  CascadeMux t734 (
    .I(net_84734),
    .O(net_84734_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b00)
  ) t736 (
    .carryinitin(),
    .carryinitout(t735)
  );
  CascadeMux t737 (
    .I(net_84839),
    .O(net_84839_cascademuxed)
  );
  CascadeMux t738 (
    .I(net_84845),
    .O(net_84845_cascademuxed)
  );
  CascadeMux t739 (
    .I(net_84851),
    .O(net_84851_cascademuxed)
  );
  CascadeMux t74 (
    .I(net_34961),
    .O(net_34961_cascademuxed)
  );
  CascadeMux t740 (
    .I(net_84863),
    .O(net_84863_cascademuxed)
  );
  CascadeMux t741 (
    .I(net_84875),
    .O(net_84875_cascademuxed)
  );
  CascadeMux t742 (
    .I(net_84980),
    .O(net_84980_cascademuxed)
  );
  CascadeMux t743 (
    .I(net_84992),
    .O(net_84992_cascademuxed)
  );
  CascadeMux t744 (
    .I(net_85004),
    .O(net_85004_cascademuxed)
  );
  CascadeMux t745 (
    .I(net_85103),
    .O(net_85103_cascademuxed)
  );
  CascadeMux t746 (
    .I(net_87692),
    .O(net_87692_cascademuxed)
  );
  CascadeMux t747 (
    .I(net_88190),
    .O(net_88190_cascademuxed)
  );
  CascadeMux t748 (
    .I(net_88208),
    .O(net_88208_cascademuxed)
  );
  CascadeMux t749 (
    .I(net_88319),
    .O(net_88319_cascademuxed)
  );
  CascadeMux t75 (
    .I(net_35060),
    .O(net_35060_cascademuxed)
  );
  CascadeMux t750 (
    .I(net_88670),
    .O(net_88670_cascademuxed)
  );
  CascadeMux t751 (
    .I(net_88676),
    .O(net_88676_cascademuxed)
  );
  CascadeMux t752 (
    .I(net_88712),
    .O(net_88712_cascademuxed)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t754 (
    .carryinitin(),
    .carryinitout(t753)
  );
  CascadeMux t756 (
    .I(net_91529),
    .O(net_91529_cascademuxed)
  );
  LocalMux t757 (
    .I(seg_2_8_lutff_2_out_7745),
    .O(seg_2_8_local_g3_2_12198)
  );
  LocalMux t758 (
    .I(seg_2_8_lutff_3_out_7746),
    .O(seg_2_8_local_g2_3_12191)
  );
  LocalMux t759 (
    .I(seg_2_8_lutff_4_out_7747),
    .O(seg_2_8_local_g2_4_12192)
  );
  CascadeMux t76 (
    .I(net_35699),
    .O(net_35699_cascademuxed)
  );
  LocalMux t760 (
    .I(seg_2_8_lutff_5_out_7748),
    .O(seg_2_8_local_g3_5_12201)
  );
  LocalMux t761 (
    .I(seg_2_8_lutff_6_out_7749),
    .O(seg_2_8_local_g0_6_12178)
  );
  LocalMux t762 (
    .I(seg_2_8_sp4_r_v_b_5_11913),
    .O(seg_2_8_local_g1_5_12185)
  );
  Span4Mux_v4 t763 (
    .I(seg_3_8_sp4_h_l_46_1816),
    .O(seg_2_8_sp4_r_v_b_5_11913)
  );
  LocalMux t764 (
    .I(seg_3_7_sp4_v_b_13_11910),
    .O(seg_3_7_local_g1_5_15893)
  );
  Span4Mux_v4 t765 (
    .I(seg_3_8_sp4_h_r_7_16106),
    .O(seg_3_7_sp4_v_b_13_11910)
  );
  Span4Mux_h4 t766 (
    .I(seg_3_8_sp4_h_l_46_1816),
    .O(seg_3_8_sp4_h_r_7_16106)
  );
  LocalMux t767 (
    .I(seg_3_8_sp4_v_b_5_11913),
    .O(seg_3_8_local_g1_5_16016)
  );
  Span4Mux_v4 t768 (
    .I(seg_3_8_sp4_h_l_46_1816),
    .O(seg_3_8_sp4_v_b_5_11913)
  );
  LocalMux t769 (
    .I(seg_5_5_sp4_h_r_31_15737),
    .O(seg_5_5_local_g3_7_23327)
  );
  CascadeMux t77 (
    .I(net_36665),
    .O(net_36665_cascademuxed)
  );
  Span4Mux_h4 t770 (
    .I(seg_3_5_sp4_v_t_39_12035),
    .O(seg_5_5_sp4_h_r_31_15737)
  );
  LocalMux t771 (
    .I(seg_4_19_sp4_h_r_24_13619),
    .O(seg_4_19_local_g3_0_21211)
  );
  LocalMux t772 (
    .I(seg_2_8_neigh_op_bnr_7_12015),
    .O(seg_2_8_local_g0_7_12179)
  );
  LocalMux t773 (
    .I(seg_3_7_lutff_7_out_12015),
    .O(seg_3_7_local_g1_7_15895)
  );
  LocalMux t774 (
    .I(seg_3_8_sp4_v_b_19_12039),
    .O(seg_3_8_local_g1_3_16014)
  );
  LocalMux t775 (
    .I(seg_2_8_neigh_op_rgt_4_12135),
    .O(seg_2_8_local_g3_4_12200)
  );
  LocalMux t776 (
    .I(seg_3_8_lutff_4_out_12135),
    .O(seg_3_8_local_g1_4_16015)
  );
  LocalMux t777 (
    .I(seg_3_13_lutff_2_out_12748),
    .O(seg_3_13_local_g0_2_16620)
  );
  LocalMux t778 (
    .I(seg_3_13_lutff_3_out_12749),
    .O(seg_3_13_local_g3_3_16645)
  );
  LocalMux t779 (
    .I(seg_3_13_lutff_4_out_12750),
    .O(seg_3_13_local_g3_4_16646)
  );
  CascadeMux t78 (
    .I(net_36671),
    .O(net_36671_cascademuxed)
  );
  LocalMux t780 (
    .I(seg_3_13_lutff_5_out_12751),
    .O(seg_3_13_local_g3_5_16647)
  );
  LocalMux t781 (
    .I(seg_3_13_lutff_6_out_12752),
    .O(seg_3_13_local_g1_6_16632)
  );
  LocalMux t782 (
    .I(seg_3_14_sp12_v_b_13_16095),
    .O(seg_3_14_local_g3_5_16770)
  );
  LocalMux t783 (
    .I(seg_8_17_sp4_h_r_33_28350),
    .O(seg_8_17_local_g2_1_35651)
  );
  Span4Mux_h4 t784 (
    .I(seg_6_17_sp4_v_b_3_24511),
    .O(seg_8_17_sp4_h_r_33_28350)
  );
  Span4Mux_v4 t785 (
    .I(seg_6_13_sp4_h_l_38_12886),
    .O(seg_6_17_sp4_v_b_3_24511)
  );
  LocalMux t786 (
    .I(seg_3_13_sp4_r_v_b_5_16359),
    .O(seg_3_13_local_g1_5_16631)
  );
  Span4Mux_v4 t787 (
    .I(seg_4_13_sp4_h_l_46_2864),
    .O(seg_3_13_sp4_r_v_b_5_16359)
  );
  LocalMux t788 (
    .I(seg_4_13_sp4_v_b_5_16359),
    .O(seg_4_13_local_g1_5_20462)
  );
  Span4Mux_v4 t789 (
    .I(seg_4_13_sp4_h_l_46_2864),
    .O(seg_4_13_sp4_v_b_5_16359)
  );
  CascadeMux t79 (
    .I(net_36689),
    .O(net_36689_cascademuxed)
  );
  LocalMux t790 (
    .I(seg_3_13_neigh_op_top_2_12871),
    .O(seg_3_13_local_g1_2_16628)
  );
  LocalMux t791 (
    .I(seg_3_14_lutff_2_out_12871),
    .O(seg_3_14_local_g2_2_16759)
  );
  LocalMux t792 (
    .I(seg_3_18_lutff_2_out_13363),
    .O(seg_3_18_local_g2_2_17251)
  );
  LocalMux t793 (
    .I(seg_4_18_neigh_op_lft_2_13363),
    .O(seg_4_18_local_g0_2_21066)
  );
  LocalMux t794 (
    .I(seg_3_18_lutff_3_out_13364),
    .O(seg_3_18_local_g2_3_17252)
  );
  LocalMux t795 (
    .I(seg_4_18_neigh_op_lft_3_13364),
    .O(seg_4_18_local_g1_3_21075)
  );
  LocalMux t796 (
    .I(seg_3_18_lutff_4_out_13365),
    .O(seg_3_18_local_g0_4_17237)
  );
  LocalMux t797 (
    .I(seg_4_18_neigh_op_lft_4_13365),
    .O(seg_4_18_local_g1_4_21076)
  );
  LocalMux t798 (
    .I(seg_3_18_lutff_5_out_13366),
    .O(seg_3_18_local_g0_5_17238)
  );
  LocalMux t799 (
    .I(seg_4_18_neigh_op_lft_5_13366),
    .O(seg_4_18_local_g0_5_21069)
  );
  CascadeMux t80 (
    .I(net_36695),
    .O(net_36695_cascademuxed)
  );
  LocalMux t800 (
    .I(seg_3_18_lutff_6_out_13367),
    .O(seg_3_18_local_g0_6_17239)
  );
  LocalMux t801 (
    .I(seg_4_18_neigh_op_lft_6_13367),
    .O(seg_4_18_local_g0_6_21070)
  );
  LocalMux t802 (
    .I(seg_3_18_lutff_7_out_13368),
    .O(seg_3_18_local_g3_7_17264)
  );
  LocalMux t803 (
    .I(seg_4_19_neigh_op_bnl_7_13368),
    .O(seg_4_19_local_g3_7_21218)
  );
  LocalMux t804 (
    .I(seg_3_19_lutff_0_out_13484),
    .O(seg_3_19_local_g1_0_17364)
  );
  LocalMux t805 (
    .I(seg_4_19_neigh_op_lft_0_13484),
    .O(seg_4_19_local_g1_0_21195)
  );
  LocalMux t806 (
    .I(seg_3_19_lutff_1_out_13485),
    .O(seg_3_19_local_g0_1_17357)
  );
  LocalMux t807 (
    .I(seg_4_18_neigh_op_tnl_1_13485),
    .O(seg_4_18_local_g3_1_21089)
  );
  LocalMux t808 (
    .I(seg_3_19_lutff_2_out_13486),
    .O(seg_3_19_local_g3_2_17382)
  );
  LocalMux t809 (
    .I(seg_4_19_neigh_op_lft_2_13486),
    .O(seg_4_19_local_g1_2_21197)
  );
  LocalMux t810 (
    .I(seg_3_19_lutff_3_out_13487),
    .O(seg_3_19_local_g1_3_17367)
  );
  LocalMux t811 (
    .I(seg_4_19_neigh_op_lft_3_13487),
    .O(seg_4_19_local_g0_3_21190)
  );
  LocalMux t812 (
    .I(seg_2_19_neigh_op_rgt_4_13488),
    .O(seg_2_19_local_g2_4_13545)
  );
  LocalMux t813 (
    .I(seg_3_19_lutff_4_out_13488),
    .O(seg_3_19_local_g2_4_17376)
  );
  LocalMux t814 (
    .I(seg_2_19_neigh_op_rgt_5_13489),
    .O(seg_2_19_local_g3_5_13554)
  );
  LocalMux t815 (
    .I(seg_3_19_lutff_5_out_13489),
    .O(seg_3_19_local_g2_5_17377)
  );
  LocalMux t816 (
    .I(seg_2_19_neigh_op_rgt_6_13490),
    .O(seg_2_19_local_g3_6_13555)
  );
  LocalMux t817 (
    .I(seg_3_19_lutff_6_out_13490),
    .O(seg_3_19_local_g0_6_17362)
  );
  LocalMux t818 (
    .I(seg_3_19_lutff_7_out_13491),
    .O(seg_3_19_local_g2_7_17379)
  );
  LocalMux t819 (
    .I(seg_4_19_neigh_op_lft_7_13491),
    .O(seg_4_19_local_g1_7_21202)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t82 (
    .carryinitin(),
    .carryinitout(t81)
  );
  LocalMux t820 (
    .I(seg_3_20_lutff_0_out_13607),
    .O(seg_3_20_local_g2_0_17495)
  );
  LocalMux t821 (
    .I(seg_4_19_neigh_op_tnl_0_13607),
    .O(seg_4_19_local_g2_0_21203)
  );
  LocalMux t822 (
    .I(seg_3_20_lutff_1_out_13608),
    .O(seg_3_20_local_g3_1_17504)
  );
  LocalMux t823 (
    .I(seg_4_20_neigh_op_lft_1_13608),
    .O(seg_4_20_local_g1_1_21319)
  );
  LocalMux t824 (
    .I(seg_2_19_neigh_op_tnr_2_13609),
    .O(seg_2_19_local_g3_2_13551)
  );
  LocalMux t825 (
    .I(seg_3_20_lutff_2_out_13609),
    .O(seg_3_20_local_g0_2_17481)
  );
  LocalMux t826 (
    .I(seg_3_20_lutff_3_out_13610),
    .O(seg_3_20_local_g3_3_17506)
  );
  LocalMux t827 (
    .I(seg_4_20_neigh_op_lft_3_13610),
    .O(seg_4_20_local_g0_3_21313)
  );
  LocalMux t828 (
    .I(seg_3_20_lutff_4_out_13611),
    .O(seg_3_20_local_g3_4_17507)
  );
  LocalMux t829 (
    .I(seg_4_20_neigh_op_lft_4_13611),
    .O(seg_4_20_local_g1_4_21322)
  );
  LocalMux t830 (
    .I(seg_3_20_lutff_5_out_13612),
    .O(seg_3_20_local_g2_5_17500)
  );
  LocalMux t831 (
    .I(seg_4_19_neigh_op_tnl_5_13612),
    .O(seg_4_19_local_g3_5_21216)
  );
  LocalMux t832 (
    .I(seg_3_20_lutff_6_out_13613),
    .O(seg_3_20_local_g1_6_17493)
  );
  LocalMux t833 (
    .I(seg_4_20_neigh_op_lft_6_13613),
    .O(seg_4_20_local_g0_6_21316)
  );
  LocalMux t834 (
    .I(seg_3_20_lutff_7_out_13614),
    .O(seg_3_20_local_g3_7_17510)
  );
  LocalMux t835 (
    .I(seg_4_19_neigh_op_tnl_7_13614),
    .O(seg_4_19_local_g2_7_21210)
  );
  LocalMux t836 (
    .I(seg_4_12_lutff_2_out_16456),
    .O(seg_4_12_local_g3_2_20352)
  );
  LocalMux t837 (
    .I(seg_5_12_neigh_op_lft_2_16456),
    .O(seg_5_12_local_g0_2_24159)
  );
  LocalMux t838 (
    .I(seg_7_12_sp4_h_r_41_20426),
    .O(seg_7_12_local_g3_1_31213)
  );
  LocalMux t839 (
    .I(seg_3_13_neigh_op_rgt_5_16582),
    .O(seg_3_13_local_g2_5_16639)
  );
  CascadeMux t84 (
    .I(net_37655),
    .O(net_37655_cascademuxed)
  );
  LocalMux t840 (
    .I(seg_4_13_lutff_5_out_16582),
    .O(seg_4_13_local_g3_5_20478)
  );
  LocalMux t841 (
    .I(seg_3_14_sp4_r_v_b_43_16854),
    .O(seg_3_14_local_g3_3_16768)
  );
  Span4Mux_v4 t842 (
    .I(seg_4_13_sp4_v_b_10_16366),
    .O(seg_3_14_sp4_r_v_b_43_16854)
  );
  LocalMux t843 (
    .I(seg_3_18_neigh_op_bnr_1_17070),
    .O(seg_3_18_local_g1_1_17242)
  );
  LocalMux t844 (
    .I(seg_4_17_lutff_1_out_17070),
    .O(seg_4_17_local_g0_1_20942)
  );
  LocalMux t845 (
    .I(seg_4_18_neigh_op_bot_1_17070),
    .O(seg_4_18_local_g0_1_21065)
  );
  LocalMux t846 (
    .I(seg_4_18_lutff_0_out_17192),
    .O(seg_4_18_local_g1_0_21072)
  );
  LocalMux t847 (
    .I(seg_4_18_lutff_6_out_17198),
    .O(seg_4_18_local_g2_6_21086)
  );
  LocalMux t848 (
    .I(seg_3_18_neigh_op_rgt_7_17199),
    .O(seg_3_18_local_g2_7_17256)
  );
  LocalMux t849 (
    .I(seg_4_18_lutff_7_out_17199),
    .O(seg_4_18_local_g2_7_21087)
  );
  CascadeMux t85 (
    .I(net_37661),
    .O(net_37661_cascademuxed)
  );
  LocalMux t850 (
    .I(seg_16_17_sp4_v_b_17_62314),
    .O(seg_16_17_local_g0_1_66281)
  );
  Span4Mux_v4 t851 (
    .I(seg_16_18_sp4_h_l_41_51181),
    .O(seg_16_17_sp4_v_b_17_62314)
  );
  Span4Mux_h4 t852 (
    .I(seg_12_18_sp4_h_l_41_35857),
    .O(seg_16_18_sp4_h_l_41_51181)
  );
  Span4Mux_h4 t853 (
    .I(seg_8_18_sp4_h_l_41_21164),
    .O(seg_12_18_sp4_h_l_41_35857)
  );
  LocalMux t854 (
    .I(seg_21_18_sp4_h_r_14_81195),
    .O(seg_21_18_local_g1_6_84941)
  );
  Span4Mux_h4 t855 (
    .I(seg_20_18_sp4_h_l_37_66497),
    .O(seg_21_18_sp4_h_r_14_81195)
  );
  Span4Mux_h4 t856 (
    .I(seg_16_18_sp4_h_l_41_51181),
    .O(seg_20_18_sp4_h_l_37_66497)
  );
  LocalMux t857 (
    .I(seg_18_19_sp4_h_r_23_70453),
    .O(seg_18_19_local_g0_7_74195)
  );
  Span4Mux_h4 t858 (
    .I(seg_17_19_sp4_h_l_42_55138),
    .O(seg_18_19_sp4_h_r_23_70453)
  );
  Span4Mux_h4 t859 (
    .I(seg_13_19_sp4_h_l_41_39811),
    .O(seg_17_19_sp4_h_l_42_55138)
  );
  CascadeMux t86 (
    .I(net_37667),
    .O(net_37667_cascademuxed)
  );
  Span4Mux_h4 t860 (
    .I(seg_9_19_sp4_h_l_45_25122),
    .O(seg_13_19_sp4_h_l_41_39811)
  );
  Span4Mux_h4 t861 (
    .I(seg_5_19_sp4_v_b_8_20933),
    .O(seg_9_19_sp4_h_l_45_25122)
  );
  LocalMux t862 (
    .I(seg_21_19_sp4_h_r_6_85152),
    .O(seg_21_19_local_g1_6_85064)
  );
  Span4Mux_h4 t863 (
    .I(seg_21_19_sp4_h_l_47_70453),
    .O(seg_21_19_sp4_h_r_6_85152)
  );
  Span4Mux_h4 t864 (
    .I(seg_17_19_sp4_h_l_42_55138),
    .O(seg_21_19_sp4_h_l_47_70453)
  );
  LocalMux t865 (
    .I(seg_21_16_sp4_v_b_13_80711),
    .O(seg_21_16_local_g1_5_84694)
  );
  Span4Mux_v4 t866 (
    .I(seg_21_17_sp4_h_l_37_70205),
    .O(seg_21_16_sp4_v_b_13_80711)
  );
  Span4Mux_h4 t867 (
    .I(seg_17_17_sp4_h_l_44_54894),
    .O(seg_21_17_sp4_h_l_37_70205)
  );
  Span4Mux_h4 t868 (
    .I(seg_13_17_sp4_h_l_36_39560),
    .O(seg_17_17_sp4_h_l_44_54894)
  );
  Span4Mux_h4 t869 (
    .I(seg_9_17_sp4_h_l_40_24873),
    .O(seg_13_17_sp4_h_l_36_39560)
  );
  CascadeMux t87 (
    .I(net_37673),
    .O(net_37673_cascademuxed)
  );
  Span4Mux_h4 t870 (
    .I(seg_5_17_sp4_v_t_37_21171),
    .O(seg_9_17_sp4_h_l_40_24873)
  );
  GlobalMux t871 (
    .I(seg_6_0_local_g1_6_26551_i3),
    .O(seg_17_13_glb_netwk_6_11)
  );
  gio2CtrlBuf t872 (
    .I(seg_6_0_local_g1_6_26551_i2),
    .O(seg_6_0_local_g1_6_26551_i3)
  );
  ICE_GB t873 (
    .GLOBALBUFFEROUTPUT(seg_6_0_local_g1_6_26551_i2),
    .USERSIGNALTOGLOBALBUFFER(seg_6_0_local_g1_6_26551_i1)
  );
  IoInMux t874 (
    .I(seg_6_0_local_g1_6_26551),
    .O(seg_6_0_local_g1_6_26551_i1)
  );
  LocalMux t875 (
    .I(seg_6_0_span4_horz_r_6_22756),
    .O(seg_6_0_local_g1_6_26551)
  );
  IoSpan4Mux t876 (
    .I(seg_5_0_span4_vert_13_19048),
    .O(seg_6_0_span4_horz_r_6_22756)
  );
  Span4Mux_v4 t877 (
    .I(seg_5_2_sp4_v_t_44_19333),
    .O(seg_5_0_span4_vert_13_19048)
  );
  Span4Mux_v4 t878 (
    .I(seg_5_6_sp4_v_t_36_19817),
    .O(seg_5_2_sp4_v_t_44_19333)
  );
  Span4Mux_v4 t879 (
    .I(seg_5_10_sp4_v_t_40_20313),
    .O(seg_5_6_sp4_v_t_36_19817)
  );
  CascadeMux t88 (
    .I(net_37679),
    .O(net_37679_cascademuxed)
  );
  Span4Mux_v4 t880 (
    .I(seg_5_14_sp4_v_t_40_20805),
    .O(seg_5_10_sp4_v_t_40_20313)
  );
  LocalMux t881 (
    .I(seg_18_10_sp4_h_r_17_69350),
    .O(seg_18_10_local_g1_1_73090)
  );
  Span4Mux_h4 t882 (
    .I(seg_17_10_sp4_h_l_36_54023),
    .O(seg_18_10_sp4_h_r_17_69350)
  );
  Span4Mux_h4 t883 (
    .I(seg_13_10_sp4_h_l_36_38699),
    .O(seg_17_10_sp4_h_l_36_54023)
  );
  Span4Mux_h4 t884 (
    .I(seg_9_10_sp4_h_l_40_24012),
    .O(seg_13_10_sp4_h_l_36_38699)
  );
  Span4Mux_h4 t885 (
    .I(seg_5_10_sp4_v_t_40_20313),
    .O(seg_9_10_sp4_h_l_40_24012)
  );
  LocalMux t886 (
    .I(seg_20_10_sp4_h_r_41_69350),
    .O(seg_20_10_local_g2_1_80129)
  );
  Span4Mux_h4 t887 (
    .I(seg_17_10_sp4_h_l_36_54023),
    .O(seg_20_10_sp4_h_r_41_69350)
  );
  LocalMux t888 (
    .I(seg_4_17_sp4_v_b_27_17095),
    .O(seg_4_17_local_g3_3_20968)
  );
  LocalMux t889 (
    .I(seg_4_18_neigh_op_top_1_17316),
    .O(seg_4_18_local_g1_1_21073)
  );
  CascadeMux t89 (
    .I(net_37691),
    .O(net_37691_cascademuxed)
  );
  LocalMux t890 (
    .I(seg_4_19_lutff_2_out_17317),
    .O(seg_4_19_local_g0_2_21189)
  );
  LocalMux t891 (
    .I(seg_4_19_lutff_4_out_17319),
    .O(seg_4_19_local_g1_4_21199)
  );
  LocalMux t892 (
    .I(seg_4_19_neigh_op_top_1_17439),
    .O(seg_4_19_local_g1_1_21196)
  );
  LocalMux t893 (
    .I(seg_8_2_sp4_r_v_b_43_33902),
    .O(seg_8_2_local_g3_3_33816)
  );
  Span4Mux_v4 t894 (
    .I(seg_9_5_sp4_h_l_37_23390),
    .O(seg_8_2_sp4_r_v_b_43_33902)
  );
  LocalMux t895 (
    .I(seg_8_3_sp4_r_v_b_24_33896),
    .O(seg_8_3_local_g0_0_33912)
  );
  Span4Mux_v4 t896 (
    .I(seg_9_5_sp4_h_l_37_23390),
    .O(seg_8_3_sp4_r_v_b_24_33896)
  );
  LocalMux t897 (
    .I(seg_9_3_sp4_v_b_24_33896),
    .O(seg_9_3_local_g2_0_37759)
  );
  Span4Mux_v4 t898 (
    .I(seg_9_5_sp4_h_l_37_23390),
    .O(seg_9_3_sp4_v_b_24_33896)
  );
  LocalMux t899 (
    .I(seg_9_4_sp4_v_b_19_33902),
    .O(seg_9_4_local_g1_3_37877)
  );
  ICE_CARRY_IN_MUX #(
    .C_INIT(2'b01)
  ) t9 (
    .carryinitin(),
    .carryinitout(t8)
  );
  CascadeMux t90 (
    .I(net_37778),
    .O(net_37778_cascademuxed)
  );
  Span4Mux_v4 t900 (
    .I(seg_9_5_sp4_h_l_37_23390),
    .O(seg_9_4_sp4_v_b_19_33902)
  );
  LocalMux t901 (
    .I(seg_9_2_sp4_h_r_44_26820),
    .O(seg_9_2_local_g3_4_37648)
  );
  Span4Mux_h4 t902 (
    .I(seg_6_2_sp4_v_t_41_23161),
    .O(seg_9_2_sp4_h_r_44_26820)
  );
  LocalMux t903 (
    .I(seg_5_12_lutff_2_out_20287),
    .O(seg_5_12_local_g2_2_24175)
  );
  LocalMux t904 (
    .I(seg_7_12_sp4_h_r_28_24257),
    .O(seg_7_12_local_g2_4_31208)
  );
  LocalMux t905 (
    .I(seg_14_20_sp4_h_r_18_55261),
    .O(seg_14_20_local_g0_2_58990)
  );
  Span4Mux_h4 t906 (
    .I(seg_13_20_sp4_h_l_42_39937),
    .O(seg_14_20_sp4_h_r_18_55261)
  );
  Span4Mux_h4 t907 (
    .I(seg_9_20_sp4_h_l_41_25241),
    .O(seg_13_20_sp4_h_l_42_39937)
  );
  LocalMux t908 (
    .I(seg_9_10_sp12_h_r_6_27622),
    .O(seg_9_10_local_g0_6_38610)
  );
  Span12Mux_h12 t909 (
    .I(seg_6_10_sp12_v_b_1_26571),
    .O(seg_9_10_sp12_h_r_6_27622)
  );
  CascadeMux t91 (
    .I(net_37784),
    .O(net_37784_cascademuxed)
  );
  LocalMux t910 (
    .I(seg_9_10_sp4_r_v_b_23_38475),
    .O(seg_9_10_local_g3_7_38635)
  );
  Span4Mux_v4 t911 (
    .I(seg_10_7_sp4_v_b_2_37975),
    .O(seg_9_10_sp4_r_v_b_23_38475)
  );
  Span4Mux_v4 t912 (
    .I(seg_10_3_sp4_h_l_39_26915),
    .O(seg_10_7_sp4_v_b_2_37975)
  );
  Span4Mux_h4 t913 (
    .I(seg_6_3_sp4_v_b_8_22900),
    .O(seg_10_3_sp4_h_l_39_26915)
  );
  LocalMux t914 (
    .I(seg_9_11_sp4_r_v_b_10_38475),
    .O(seg_9_11_local_g2_2_38745)
  );
  Span4Mux_v4 t915 (
    .I(seg_10_7_sp4_v_b_2_37975),
    .O(seg_9_11_sp4_r_v_b_10_38475)
  );
  LocalMux t916 (
    .I(seg_8_2_sp4_h_r_16_30059),
    .O(seg_8_2_local_g1_0_33797)
  );
  Span4Mux_h4 t917 (
    .I(seg_7_2_sp4_v_b_5_26691),
    .O(seg_8_2_sp4_h_r_16_30059)
  );
  LocalMux t918 (
    .I(seg_7_12_lutff_2_out_27687),
    .O(seg_7_12_local_g3_2_31214)
  );
  LocalMux t919 (
    .I(seg_7_12_lutff_3_out_27688),
    .O(seg_7_12_local_g2_3_31207)
  );
  CascadeMux t92 (
    .I(net_37790),
    .O(net_37790_cascademuxed)
  );
  LocalMux t920 (
    .I(seg_9_12_sp4_h_r_34_31284),
    .O(seg_9_12_local_g2_2_38868)
  );
  LocalMux t921 (
    .I(seg_9_3_neigh_op_bnl_1_29882),
    .O(seg_9_3_local_g3_1_37768)
  );
  LocalMux t922 (
    .I(seg_8_2_lutff_2_out_29883),
    .O(seg_8_2_local_g0_2_33791)
  );
  LocalMux t923 (
    .I(seg_7_1_neigh_op_tnr_3_29884),
    .O(seg_7_1_local_g2_3_29814)
  );
  LocalMux t924 (
    .I(seg_9_2_neigh_op_lft_3_29884),
    .O(seg_9_2_local_g0_3_37623)
  );
  LocalMux t925 (
    .I(seg_8_2_lutff_6_out_29887),
    .O(seg_8_2_local_g1_6_33803)
  );
  LocalMux t926 (
    .I(seg_7_1_neigh_op_tnr_7_29888),
    .O(seg_7_1_local_g3_7_29826)
  );
  LocalMux t927 (
    .I(seg_6_0_span4_vert_18_22884),
    .O(seg_6_0_local_g0_2_26539)
  );
  Span4Mux_v4 t928 (
    .I(seg_6_2_sp4_h_r_2_26813),
    .O(seg_6_0_span4_vert_18_22884)
  );
  LocalMux t929 (
    .I(seg_7_0_span4_horz_r_14_18925),
    .O(seg_7_0_local_g0_6_29743)
  );
  CascadeMux t93 (
    .I(net_37796),
    .O(net_37796_cascademuxed)
  );
  IoSpan4Mux t930 (
    .I(seg_8_0_span4_vert_37_29936),
    .O(seg_7_0_span4_horz_r_14_18925)
  );
  LocalMux t931 (
    .I(seg_8_3_lutff_4_out_30044),
    .O(seg_8_3_local_g0_4_33916)
  );
  LocalMux t932 (
    .I(seg_8_2_neigh_op_top_5_30045),
    .O(seg_8_2_local_g1_5_33802)
  );
  LocalMux t933 (
    .I(seg_8_3_lutff_5_out_30045),
    .O(seg_8_3_local_g3_5_33941)
  );
  LocalMux t934 (
    .I(seg_9_2_neigh_op_tnl_5_30045),
    .O(seg_9_2_local_g3_5_37649)
  );
  LocalMux t935 (
    .I(seg_9_3_neigh_op_lft_5_30045),
    .O(seg_9_3_local_g0_5_37748)
  );
  LocalMux t936 (
    .I(seg_9_4_neigh_op_bnl_5_30045),
    .O(seg_9_4_local_g3_5_37895)
  );
  LocalMux t937 (
    .I(seg_8_3_lutff_6_out_30046),
    .O(seg_8_3_local_g1_6_33926)
  );
  LocalMux t938 (
    .I(seg_8_3_sp4_h_r_18_30184),
    .O(seg_8_3_local_g0_2_33914)
  );
  LocalMux t939 (
    .I(seg_10_2_sp4_v_b_19_37591),
    .O(seg_10_2_local_g1_3_41462)
  );
  CascadeMux t94 (
    .I(net_37802),
    .O(net_37802_cascademuxed)
  );
  Span4Mux_v4 t940 (
    .I(seg_10_3_sp4_h_l_43_26919),
    .O(seg_10_2_sp4_v_b_19_37591)
  );
  LocalMux t941 (
    .I(seg_10_3_sp4_h_r_2_41672),
    .O(seg_10_3_local_g0_2_41576)
  );
  Span4Mux_h4 t942 (
    .I(seg_10_3_sp4_h_l_43_26919),
    .O(seg_10_3_sp4_h_r_2_41672)
  );
  LocalMux t943 (
    .I(seg_9_3_sp4_v_b_19_33774),
    .O(seg_9_3_local_g1_3_37754)
  );
  LocalMux t944 (
    .I(seg_9_5_neigh_op_bnl_1_30164),
    .O(seg_9_5_local_g3_1_38014)
  );
  LocalMux t945 (
    .I(seg_8_12_sp12_v_b_2_33722),
    .O(seg_8_12_local_g3_2_35045)
  );
  LocalMux t946 (
    .I(seg_8_23_sp12_v_b_5_35234),
    .O(seg_8_23_local_g2_5_36393)
  );
  Span12Mux_v12 t947 (
    .I(seg_8_13_sp12_v_b_1_33722),
    .O(seg_8_23_sp12_v_b_5_35234)
  );
  LocalMux t948 (
    .I(seg_8_31_span12_vert_13_36710),
    .O(seg_8_31_local_g1_5_37382)
  );
  Span12Mux_v12 t949 (
    .I(seg_8_25_sp12_v_b_1_35234),
    .O(seg_8_31_span12_vert_13_36710)
  );
  CascadeMux t95 (
    .I(net_37808),
    .O(net_37808_cascademuxed)
  );
  Span12Mux_v12 t950 (
    .I(seg_8_13_sp12_v_b_1_33722),
    .O(seg_8_25_sp12_v_b_1_35234)
  );
  LocalMux t951 (
    .I(seg_9_28_sp4_h_r_16_37088),
    .O(seg_9_28_local_g0_0_40818)
  );
  Span4Mux_h4 t952 (
    .I(seg_8_28_sp4_v_b_11_32903),
    .O(seg_9_28_sp4_h_r_16_37088)
  );
  Span4Mux_v4 t953 (
    .I(seg_8_24_sp4_v_b_3_32403),
    .O(seg_8_28_sp4_v_b_11_32903)
  );
  Sp12to4 t954 (
    .I(seg_8_23_sp12_v_b_5_35234),
    .O(seg_8_24_sp4_v_b_3_32403)
  );
  LocalMux t955 (
    .I(seg_9_28_sp4_h_r_16_37088),
    .O(seg_9_28_local_g1_0_40826)
  );
  LocalMux t956 (
    .I(seg_15_25_sp12_h_r_14_36709),
    .O(seg_15_25_local_g0_6_63439)
  );
  Span12Mux_h12 t957 (
    .I(seg_8_25_sp12_v_b_1_35234),
    .O(seg_15_25_sp12_h_r_14_36709)
  );
  LocalMux t958 (
    .I(seg_18_31_span4_vert_34_71823),
    .O(seg_18_31_local_g0_2_75679)
  );
  Span4Mux_v4 t959 (
    .I(seg_18_29_sp4_v_b_10_71335),
    .O(seg_18_31_span4_vert_34_71823)
  );
  CascadeMux t96 (
    .I(net_37814),
    .O(net_37814_cascademuxed)
  );
  Span4Mux_v4 t960 (
    .I(seg_18_25_sp4_h_r_10_75022),
    .O(seg_18_29_sp4_v_b_10_71335)
  );
  Sp12to4 t961 (
    .I(seg_19_25_sp12_h_r_22_36709),
    .O(seg_18_25_sp4_h_r_10_75022)
  );
  Span12Mux_h12 t962 (
    .I(seg_8_25_sp12_v_b_1_35234),
    .O(seg_19_25_sp12_h_r_22_36709)
  );
  LocalMux t963 (
    .I(seg_3_7_sp4_v_b_23_11920),
    .O(seg_3_7_local_g0_7_15887)
  );
  Span4Mux_v4 t964 (
    .I(seg_3_4_sp4_h_r_10_15607),
    .O(seg_3_7_sp4_v_b_23_11920)
  );
  Span4Mux_h4 t965 (
    .I(seg_7_4_sp4_h_r_7_30307),
    .O(seg_3_4_sp4_h_r_10_15607)
  );
  LocalMux t966 (
    .I(seg_4_12_sp4_h_r_15_16593),
    .O(seg_4_12_local_g1_7_20341)
  );
  Span4Mux_h4 t967 (
    .I(seg_7_12_sp4_v_b_9_27543),
    .O(seg_4_12_sp4_h_r_15_16593)
  );
  Span4Mux_v4 t968 (
    .I(seg_7_8_sp4_v_b_1_27127),
    .O(seg_7_12_sp4_v_b_9_27543)
  );
  Span4Mux_v4 t969 (
    .I(seg_7_4_sp4_h_r_7_30307),
    .O(seg_7_8_sp4_v_b_1_27127)
  );
  CascadeMux t97 (
    .I(net_37820),
    .O(net_37820_cascademuxed)
  );
  LocalMux t970 (
    .I(seg_7_0_span4_vert_42_26720),
    .O(seg_7_0_local_g1_2_29747)
  );
  Span4Mux_v4 t971 (
    .I(seg_7_4_sp4_h_r_7_30307),
    .O(seg_7_0_span4_vert_42_26720)
  );
  LocalMux t972 (
    .I(seg_10_3_sp4_r_v_b_18_41435),
    .O(seg_10_3_local_g3_2_41600)
  );
  Span4Mux_v4 t973 (
    .I(seg_11_4_sp4_h_l_42_30307),
    .O(seg_10_3_sp4_r_v_b_18_41435)
  );
  LocalMux t974 (
    .I(seg_10_11_sp4_r_v_b_21_42427),
    .O(seg_10_11_local_g3_5_42587)
  );
  Span4Mux_v4 t975 (
    .I(seg_11_8_sp4_v_b_0_41927),
    .O(seg_10_11_sp4_r_v_b_21_42427)
  );
  Span4Mux_v4 t976 (
    .I(seg_11_4_sp4_h_l_42_30307),
    .O(seg_11_8_sp4_v_b_0_41927)
  );
  LocalMux t977 (
    .I(seg_14_3_sp4_r_v_b_12_56751),
    .O(seg_14_3_local_g2_4_56917)
  );
  Span4Mux_v4 t978 (
    .I(seg_15_4_sp4_h_l_42_45631),
    .O(seg_14_3_sp4_r_v_b_12_56751)
  );
  Span4Mux_h4 t979 (
    .I(seg_11_4_sp4_h_l_42_30307),
    .O(seg_15_4_sp4_h_l_42_45631)
  );
  CascadeMux t98 (
    .I(net_37901),
    .O(net_37901_cascademuxed)
  );
  LocalMux t980 (
    .I(seg_14_7_sp4_r_v_b_18_57255),
    .O(seg_14_7_local_g3_2_57415)
  );
  Span4Mux_v4 t981 (
    .I(seg_15_4_sp4_h_l_42_45631),
    .O(seg_14_7_sp4_r_v_b_18_57255)
  );
  LocalMux t982 (
    .I(seg_15_6_sp4_v_b_31_57255),
    .O(seg_15_6_local_g2_7_61119)
  );
  Span4Mux_v4 t983 (
    .I(seg_15_4_sp4_h_l_42_45631),
    .O(seg_15_6_sp4_v_b_31_57255)
  );
  LocalMux t984 (
    .I(seg_19_14_sp4_v_b_35_73566),
    .O(seg_19_14_local_g3_3_77156)
  );
  Span4Mux_v4 t985 (
    .I(seg_19_12_sp4_v_b_11_73074),
    .O(seg_19_14_sp4_v_b_35_73566)
  );
  Span4Mux_v4 t986 (
    .I(seg_19_8_sp4_v_b_3_72574),
    .O(seg_19_12_sp4_v_b_11_73074)
  );
  Span4Mux_v4 t987 (
    .I(seg_19_4_sp4_h_l_47_60946),
    .O(seg_19_8_sp4_v_b_3_72574)
  );
  Span4Mux_h4 t988 (
    .I(seg_15_4_sp4_h_l_42_45631),
    .O(seg_19_4_sp4_h_l_47_60946)
  );
  LocalMux t989 (
    .I(seg_19_15_sp4_v_b_18_73562),
    .O(seg_19_15_local_g0_2_77233)
  );
  CascadeMux t99 (
    .I(net_37931),
    .O(net_37931_cascademuxed)
  );
  Span4Mux_v4 t990 (
    .I(seg_19_12_sp4_v_b_11_73074),
    .O(seg_19_15_sp4_v_b_18_73562)
  );
  LocalMux t991 (
    .I(seg_19_15_sp4_v_b_20_73564),
    .O(seg_19_15_local_g0_4_77235)
  );
  Span4Mux_v4 t992 (
    .I(seg_19_12_sp4_v_b_6_73071),
    .O(seg_19_15_sp4_v_b_20_73564)
  );
  Span4Mux_v4 t993 (
    .I(seg_19_8_sp4_v_b_3_72574),
    .O(seg_19_12_sp4_v_b_6_73071)
  );
  LocalMux t994 (
    .I(seg_11_7_sp4_r_v_b_18_45763),
    .O(seg_11_7_local_g3_2_45923)
  );
  Span4Mux_v4 t995 (
    .I(seg_12_4_sp4_h_l_39_34133),
    .O(seg_11_7_sp4_r_v_b_18_45763)
  );
  LocalMux t996 (
    .I(seg_11_8_sp4_r_v_b_2_45760),
    .O(seg_11_8_local_g1_2_46030)
  );
  Span4Mux_v4 t997 (
    .I(seg_12_4_sp4_h_l_39_34133),
    .O(seg_11_8_sp4_r_v_b_2_45760)
  );
  LocalMux t998 (
    .I(seg_11_8_sp4_r_v_b_7_45763),
    .O(seg_11_8_local_g1_7_46035)
  );
  Span4Mux_v4 t999 (
    .I(seg_12_4_sp4_h_l_39_34133),
    .O(seg_11_8_sp4_r_v_b_7_45763)
  );
endmodule
