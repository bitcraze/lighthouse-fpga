/* verilator lint_off UNUSED */
/* verilator lint_off UNDRIVEN */
(* blackbox, keep *)
module SB_WARMBOOT (
	input BOOT,
	input S1,
	input S0
);
endmodule
/* verilator lint_on UNUSED */
/* verilator lint_on UNDRIVEN */
